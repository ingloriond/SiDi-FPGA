
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity basic is
port(
        clock:in std_logic;
	we:in std_logic;
        data:in std_logic_vector(7 downto 0);
        address:in std_logic_vector(12 downto 0);
        q:out std_logic_vector(7 downto 0)
);
end basic;

architecture syn of basic is
        type rom_type is array(0 to 8191) of std_logic_vector(7 downto 0);
        signal ROM:rom_type:=
(
	X"a5",
X"ca",
X"d0",
X"04",
X"a5",
X"08",
X"d0",
X"45",
X"a2",
X"ff",
X"9a",
X"d8",
X"ae",
X"e7",
X"02",
X"ac",
X"e8",
X"02",
X"86",
X"80",
X"84",
X"81",
X"a9",
X"00",
X"85",
X"92",
X"85",
X"ca",
X"c8",
X"8a",
X"a2",
X"82",
X"95",
X"00",
X"e8",
X"94",
X"00",
X"e8",
X"e0",
X"92",
X"90",
X"f6",
X"a2",
X"86",
X"a0",
X"01",
X"20",
X"7a",
X"a8",
X"a2",
X"8c",
X"a0",
X"03",
X"20",
X"7a",
X"a8",
X"a9",
X"00",
X"a8",
X"91",
X"84",
X"91",
X"8a",
X"c8",
X"a9",
X"80",
X"91",
X"8a",
X"c8",
X"a9",
X"03",
X"91",
X"8a",
X"a9",
X"0a",
X"85",
X"c9",
X"20",
X"f1",
X"b8",
X"20",
X"45",
X"bd",
X"20",
X"5b",
X"bd",
X"a5",
X"92",
X"f0",
X"03",
X"20",
X"9d",
X"bd",
X"20",
X"62",
X"bd",
X"a5",
X"ca",
X"d0",
X"9c",
X"a2",
X"ff",
X"9a",
X"20",
X"51",
X"da",
X"a9",
X"5d",
X"85",
X"c2",
X"20",
X"ed",
X"bd",
X"20",
X"f2",
X"a9",
X"f0",
X"ea",
X"a9",
X"00",
X"85",
X"f2",
X"85",
X"9f",
X"85",
X"94",
X"85",
X"a6",
X"85",
X"b3",
X"85",
X"b0",
X"85",
X"b1",
X"a5",
X"84",
X"85",
X"ad",
X"a5",
X"85",
X"85",
X"ae",
X"20",
X"a1",
X"db",
X"20",
X"9a",
X"a1",
X"20",
X"c4",
X"a2",
X"a5",
X"d5",
X"10",
X"02",
X"85",
X"a6",
X"20",
X"a1",
X"db",
X"a4",
X"f2",
X"84",
X"a8",
X"b1",
X"f3",
X"c9",
X"9b",
X"d0",
X"07",
X"24",
X"a6",
X"30",
X"b2",
X"4c",
X"86",
X"a1",
X"a5",
X"94",
X"85",
X"a7",
X"20",
X"c4",
X"a2",
X"20",
X"a1",
X"db",
X"a9",
X"a4",
X"a0",
X"9f",
X"a2",
X"02",
X"20",
X"54",
X"a4",
X"86",
X"f2",
X"a5",
X"af",
X"20",
X"c4",
X"a2",
X"20",
X"a1",
X"db",
X"20",
X"be",
X"a1",
X"90",
X"35",
X"a4",
X"9f",
X"b1",
X"f3",
X"c9",
X"9b",
X"d0",
X"06",
X"c8",
X"91",
X"f3",
X"88",
X"a9",
X"20",
X"09",
X"80",
X"91",
X"f3",
X"a9",
X"40",
X"05",
X"a6",
X"85",
X"a6",
X"a4",
X"a8",
X"84",
X"f2",
X"a2",
X"03",
X"86",
X"a7",
X"e8",
X"86",
X"94",
X"a9",
X"37",
X"20",
X"c4",
X"a2",
X"a4",
X"f2",
X"b1",
X"f3",
X"e6",
X"f2",
X"c9",
X"9b",
X"d0",
X"f3",
X"20",
X"c4",
X"a2",
X"a5",
X"94",
X"a4",
X"a7",
X"91",
X"80",
X"a4",
X"f2",
X"88",
X"b1",
X"f3",
X"c9",
X"9b",
X"d0",
X"9a",
X"a0",
X"02",
X"a5",
X"94",
X"91",
X"80",
X"20",
X"a2",
X"a9",
X"a9",
X"00",
X"b0",
X"03",
X"20",
X"dc",
X"a9",
X"38",
X"e5",
X"94",
X"f0",
X"1e",
X"b0",
X"13",
X"49",
X"ff",
X"a8",
X"c8",
X"a2",
X"8a",
X"20",
X"7a",
X"a8",
X"a5",
X"97",
X"85",
X"8a",
X"a5",
X"98",
X"85",
X"8b",
X"d0",
X"09",
X"a8",
X"20",
X"d0",
X"a9",
X"a2",
X"8a",
X"20",
X"f8",
X"a8",
X"a4",
X"94",
X"88",
X"b1",
X"80",
X"91",
X"8a",
X"98",
X"d0",
X"f8",
X"24",
X"a6",
X"50",
X"29",
X"a5",
X"b1",
X"0a",
X"0a",
X"0a",
X"a2",
X"88",
X"20",
X"f7",
X"a8",
X"38",
X"a5",
X"84",
X"e5",
X"ad",
X"a8",
X"a5",
X"85",
X"e5",
X"ae",
X"a2",
X"84",
X"20",
X"fa",
X"a8",
X"24",
X"a6",
X"10",
X"06",
X"20",
X"aa",
X"b5",
X"4c",
X"60",
X"a0",
X"20",
X"8e",
X"b5",
X"4c",
X"60",
X"a0",
X"10",
X"fb",
X"4c",
X"5e",
X"a9",
X"20",
X"a2",
X"a9",
X"b0",
X"f3",
X"20",
X"dc",
X"a9",
X"a8",
X"20",
X"d0",
X"a9",
X"a2",
X"8a",
X"20",
X"f8",
X"a8",
X"4c",
X"60",
X"a0",
X"20",
X"00",
X"d8",
X"90",
X"08",
X"a9",
X"00",
X"85",
X"f2",
X"a0",
X"80",
X"30",
X"09",
X"20",
X"41",
X"ad",
X"a4",
X"d5",
X"30",
X"f1",
X"a5",
X"d4",
X"84",
X"a1",
X"85",
X"a0",
X"20",
X"c4",
X"a2",
X"a5",
X"a1",
X"85",
X"d5",
X"4c",
X"c4",
X"a2",
X"a0",
X"01",
X"b1",
X"95",
X"85",
X"9e",
X"8d",
X"83",
X"04",
X"88",
X"b1",
X"95",
X"85",
X"9d",
X"8d",
X"82",
X"04",
X"84",
X"a9",
X"a5",
X"94",
X"8d",
X"81",
X"04",
X"a5",
X"f2",
X"8d",
X"80",
X"04",
X"20",
X"93",
X"a2",
X"30",
X"16",
X"c9",
X"01",
X"90",
X"24",
X"d0",
X"06",
X"20",
X"08",
X"a2",
X"4c",
X"59",
X"a2",
X"c9",
X"05",
X"90",
X"55",
X"20",
X"9b",
X"a2",
X"4c",
X"59",
X"a2",
X"38",
X"e9",
X"c1",
X"b0",
X"02",
X"a2",
X"ff",
X"18",
X"65",
X"9d",
X"48",
X"8a",
X"65",
X"9e",
X"48",
X"4c",
X"1b",
X"a2",
X"20",
X"93",
X"a2",
X"48",
X"20",
X"93",
X"a2",
X"48",
X"90",
X"09",
X"68",
X"a8",
X"68",
X"aa",
X"98",
X"48",
X"8a",
X"48",
X"60",
X"a6",
X"a9",
X"e8",
X"e8",
X"e8",
X"e8",
X"f0",
X"1f",
X"86",
X"a9",
X"a5",
X"f2",
X"9d",
X"80",
X"04",
X"a5",
X"94",
X"9d",
X"81",
X"04",
X"a5",
X"9d",
X"9d",
X"82",
X"04",
X"a5",
X"9e",
X"9d",
X"83",
X"04",
X"68",
X"85",
X"9e",
X"68",
X"85",
X"9d",
X"4c",
X"db",
X"a1",
X"4c",
X"18",
X"b9",
X"a6",
X"a9",
X"f0",
X"d1",
X"bd",
X"82",
X"04",
X"85",
X"9d",
X"bd",
X"83",
X"04",
X"85",
X"9e",
X"ca",
X"ca",
X"ca",
X"ca",
X"86",
X"a9",
X"b0",
X"03",
X"4c",
X"db",
X"a1",
X"20",
X"93",
X"a2",
X"30",
X"fb",
X"c9",
X"02",
X"b0",
X"08",
X"20",
X"8c",
X"a2",
X"20",
X"8c",
X"a2",
X"d0",
X"ef",
X"c9",
X"03",
X"f0",
X"d2",
X"b0",
X"e9",
X"a5",
X"f2",
X"c5",
X"9f",
X"90",
X"02",
X"85",
X"9f",
X"a6",
X"a9",
X"bd",
X"80",
X"04",
X"85",
X"f2",
X"bd",
X"81",
X"04",
X"85",
X"94",
X"4c",
X"db",
X"a1",
X"e6",
X"9d",
X"d0",
X"02",
X"e6",
X"9e",
X"60",
X"20",
X"8c",
X"a2",
X"a2",
X"00",
X"a1",
X"9d",
X"60",
X"c9",
X"0f",
X"f0",
X"17",
X"b0",
X"40",
X"c9",
X"0d",
X"d0",
X"06",
X"20",
X"8c",
X"a2",
X"4c",
X"e4",
X"a2",
X"68",
X"68",
X"a9",
X"04",
X"48",
X"a9",
X"a6",
X"48",
X"4c",
X"1b",
X"a2",
X"20",
X"8c",
X"a2",
X"a0",
X"00",
X"b1",
X"9d",
X"a4",
X"94",
X"88",
X"91",
X"80",
X"18",
X"60",
X"a4",
X"94",
X"91",
X"80",
X"e6",
X"94",
X"d0",
X"f7",
X"4c",
X"18",
X"b9",
X"a2",
X"ff",
X"9a",
X"a5",
X"94",
X"a4",
X"a7",
X"91",
X"80",
X"4c",
X"b1",
X"a0",
X"a2",
X"ff",
X"9a",
X"4c",
X"fb",
X"a0",
X"20",
X"a1",
X"db",
X"a5",
X"f2",
X"c5",
X"b3",
X"f0",
X"15",
X"85",
X"b3",
X"a9",
X"a7",
X"a0",
X"de",
X"a2",
X"00",
X"20",
X"54",
X"a4",
X"b0",
X"23",
X"86",
X"b2",
X"a5",
X"af",
X"69",
X"10",
X"85",
X"b0",
X"a0",
X"00",
X"b1",
X"9d",
X"c5",
X"b0",
X"f0",
X"0a",
X"c9",
X"44",
X"d0",
X"13",
X"a5",
X"b0",
X"c9",
X"44",
X"90",
X"0d",
X"20",
X"c4",
X"a2",
X"a6",
X"b2",
X"86",
X"f2",
X"18",
X"60",
X"a9",
X"00",
X"85",
X"b0",
X"38",
X"60",
X"a9",
X"00",
X"f0",
X"02",
X"a9",
X"80",
X"85",
X"d2",
X"20",
X"a1",
X"db",
X"a5",
X"f2",
X"85",
X"ac",
X"20",
X"e8",
X"a3",
X"b0",
X"25",
X"20",
X"e1",
X"a2",
X"a5",
X"b0",
X"f0",
X"08",
X"a4",
X"b2",
X"b1",
X"f3",
X"c9",
X"30",
X"90",
X"16",
X"e6",
X"f2",
X"20",
X"e8",
X"a3",
X"90",
X"f9",
X"20",
X"af",
X"db",
X"90",
X"f4",
X"b1",
X"f3",
X"c9",
X"24",
X"f0",
X"06",
X"24",
X"d2",
X"10",
X"09",
X"38",
X"60",
X"24",
X"d2",
X"10",
X"fa",
X"c8",
X"d0",
X"0d",
X"b1",
X"f3",
X"c9",
X"28",
X"d0",
X"07",
X"c8",
X"a9",
X"40",
X"05",
X"d2",
X"85",
X"d2",
X"a5",
X"ac",
X"85",
X"f2",
X"84",
X"ac",
X"a5",
X"83",
X"a4",
X"82",
X"a2",
X"00",
X"20",
X"54",
X"a4",
X"b0",
X"0a",
X"e4",
X"ac",
X"f0",
X"4d",
X"20",
X"82",
X"a4",
X"4c",
X"7e",
X"a3",
X"38",
X"a5",
X"ac",
X"e5",
X"f2",
X"85",
X"f2",
X"a8",
X"a2",
X"84",
X"20",
X"7a",
X"a8",
X"a5",
X"af",
X"85",
X"d3",
X"a4",
X"f2",
X"88",
X"a6",
X"ac",
X"ca",
X"bd",
X"80",
X"05",
X"91",
X"97",
X"ca",
X"88",
X"10",
X"f7",
X"a4",
X"f2",
X"88",
X"b1",
X"97",
X"09",
X"80",
X"91",
X"97",
X"a0",
X"08",
X"a2",
X"88",
X"20",
X"7a",
X"a8",
X"e6",
X"b1",
X"a0",
X"02",
X"a9",
X"00",
X"99",
X"d2",
X"00",
X"c8",
X"c0",
X"08",
X"90",
X"f8",
X"88",
X"b9",
X"d2",
X"00",
X"91",
X"97",
X"88",
X"10",
X"f8",
X"24",
X"d2",
X"50",
X"02",
X"c6",
X"ac",
X"a5",
X"ac",
X"85",
X"f2",
X"a5",
X"af",
X"30",
X"06",
X"09",
X"80",
X"18",
X"4c",
X"c4",
X"a2",
X"4c",
X"2c",
X"b9",
X"a4",
X"f2",
X"b1",
X"f3",
X"c9",
X"41",
X"90",
X"03",
X"c9",
X"5b",
X"60",
X"38",
X"60",
X"20",
X"a1",
X"db",
X"a5",
X"f2",
X"85",
X"ac",
X"20",
X"00",
X"d8",
X"90",
X"05",
X"a5",
X"ac",
X"85",
X"f2",
X"60",
X"a9",
X"0e",
X"20",
X"c4",
X"a2",
X"c8",
X"a2",
X"00",
X"b5",
X"d4",
X"91",
X"80",
X"c8",
X"e8",
X"e0",
X"06",
X"90",
X"f6",
X"84",
X"94",
X"18",
X"60",
X"20",
X"a1",
X"db",
X"a4",
X"f2",
X"b1",
X"f3",
X"c9",
X"22",
X"d0",
X"cc",
X"a9",
X"0f",
X"20",
X"c4",
X"a2",
X"a5",
X"94",
X"85",
X"ab",
X"20",
X"c4",
X"a2",
X"e6",
X"f2",
X"a4",
X"f2",
X"b1",
X"f3",
X"c9",
X"9b",
X"f0",
X"0c",
X"c9",
X"22",
X"f0",
X"06",
X"20",
X"c4",
X"a2",
X"4c",
X"33",
X"a4",
X"e6",
X"f2",
X"18",
X"a5",
X"94",
X"e5",
X"ab",
X"a4",
X"ab",
X"91",
X"80",
X"18",
X"60",
X"86",
X"aa",
X"a2",
X"ff",
X"86",
X"af",
X"85",
X"96",
X"84",
X"95",
X"e6",
X"af",
X"a6",
X"f2",
X"a4",
X"aa",
X"b1",
X"95",
X"f0",
X"25",
X"a9",
X"00",
X"08",
X"bd",
X"80",
X"05",
X"29",
X"7f",
X"c9",
X"2e",
X"f0",
X"1b",
X"51",
X"95",
X"0a",
X"f0",
X"02",
X"68",
X"08",
X"c8",
X"e8",
X"90",
X"ec",
X"28",
X"f0",
X"d0",
X"18",
X"98",
X"65",
X"95",
X"a8",
X"a5",
X"96",
X"69",
X"00",
X"d0",
X"cd",
X"38",
X"60",
X"a9",
X"02",
X"c5",
X"aa",
X"d0",
X"df",
X"b1",
X"95",
X"30",
X"03",
X"c8",
X"d0",
X"f9",
X"38",
X"b0",
X"dc",
X"c2",
X"a7",
X"52",
X"45",
X"cd",
X"c5",
X"a7",
X"44",
X"41",
X"54",
X"c1",
X"ee",
X"a6",
X"49",
X"4e",
X"50",
X"55",
X"d4",
X"b7",
X"a6",
X"43",
X"4f",
X"4c",
X"4f",
X"d2",
X"2c",
X"a7",
X"4c",
X"49",
X"53",
X"d4",
X"1d",
X"a7",
X"45",
X"4e",
X"54",
X"45",
X"d2",
X"ba",
X"a6",
X"4c",
X"45",
X"d4",
X"8e",
X"a7",
X"49",
X"c6",
X"cc",
X"a6",
X"46",
X"4f",
X"d2",
X"e4",
X"a6",
X"4e",
X"45",
X"58",
X"d4",
X"b7",
X"a6",
X"47",
X"4f",
X"54",
X"cf",
X"b7",
X"a6",
X"47",
X"4f",
X"20",
X"54",
X"cf",
X"b7",
X"a6",
X"47",
X"4f",
X"53",
X"55",
X"c2",
X"b7",
X"a6",
X"54",
X"52",
X"41",
X"d0",
X"b8",
X"a6",
X"42",
X"59",
X"c5",
X"b8",
X"a6",
X"43",
X"4f",
X"4e",
X"d4",
X"59",
X"a7",
X"43",
X"4f",
X"cd",
X"1a",
X"a7",
X"43",
X"4c",
X"4f",
X"53",
X"c5",
X"b8",
X"a6",
X"43",
X"4c",
X"d2",
X"b8",
X"a6",
X"44",
X"45",
X"c7",
X"59",
X"a7",
X"44",
X"49",
X"cd",
X"b8",
X"a6",
X"45",
X"4e",
X"c4",
X"b8",
X"a6",
X"4e",
X"45",
X"d7",
X"13",
X"a7",
X"4f",
X"50",
X"45",
X"ce",
X"1d",
X"a7",
X"4c",
X"4f",
X"41",
X"c4",
X"1d",
X"a7",
X"53",
X"41",
X"56",
X"c5",
X"3a",
X"a7",
X"53",
X"54",
X"41",
X"54",
X"55",
X"d3",
X"43",
X"a7",
X"4e",
X"4f",
X"54",
X"c5",
X"43",
X"a7",
X"50",
X"4f",
X"49",
X"4e",
X"d4",
X"11",
X"a7",
X"58",
X"49",
X"cf",
X"5c",
X"a7",
X"4f",
X"ce",
X"56",
X"a7",
X"50",
X"4f",
X"4b",
X"c5",
X"f6",
X"a6",
X"50",
X"52",
X"49",
X"4e",
X"d4",
X"b8",
X"a6",
X"52",
X"41",
X"c4",
X"ef",
X"a6",
X"52",
X"45",
X"41",
X"c4",
X"e9",
X"a6",
X"52",
X"45",
X"53",
X"54",
X"4f",
X"52",
X"c5",
X"b8",
X"a6",
X"52",
X"45",
X"54",
X"55",
X"52",
X"ce",
X"20",
X"a7",
X"52",
X"55",
X"ce",
X"b8",
X"a6",
X"53",
X"54",
X"4f",
X"d0",
X"b8",
X"a6",
X"50",
X"4f",
X"d0",
X"f6",
X"a6",
X"bf",
X"e2",
X"a6",
X"47",
X"45",
X"d4",
X"b4",
X"a6",
X"50",
X"55",
X"d4",
X"b7",
X"a6",
X"47",
X"52",
X"41",
X"50",
X"48",
X"49",
X"43",
X"d3",
X"56",
X"a7",
X"50",
X"4c",
X"4f",
X"d4",
X"56",
X"a7",
X"50",
X"4f",
X"53",
X"49",
X"54",
X"49",
X"4f",
X"ce",
X"b8",
X"a6",
X"44",
X"4f",
X"d3",
X"56",
X"a7",
X"44",
X"52",
X"41",
X"57",
X"54",
X"cf",
X"54",
X"a7",
X"53",
X"45",
X"54",
X"43",
X"4f",
X"4c",
X"4f",
X"d2",
X"dc",
X"a6",
X"4c",
X"4f",
X"43",
X"41",
X"54",
X"c5",
X"52",
X"a7",
X"53",
X"4f",
X"55",
X"4e",
X"c4",
X"fa",
X"a6",
X"4c",
X"50",
X"52",
X"49",
X"4e",
X"d4",
X"b8",
X"a6",
X"43",
X"53",
X"41",
X"56",
X"c5",
X"b8",
X"a6",
X"43",
X"4c",
X"4f",
X"41",
X"c4",
X"ba",
X"a6",
X"00",
X"80",
X"00",
X"2a",
X"45",
X"52",
X"52",
X"4f",
X"52",
X"2d",
X"20",
X"a0",
X"53",
X"54",
X"4f",
X"50",
X"50",
X"45",
X"44",
X"a0",
X"cd",
X"c4",
X"02",
X"c2",
X"03",
X"2b",
X"ba",
X"2c",
X"db",
X"02",
X"cd",
X"d8",
X"03",
X"25",
X"0f",
X"35",
X"02",
X"26",
X"0f",
X"36",
X"02",
X"28",
X"03",
X"fe",
X"02",
X"e8",
X"02",
X"01",
X"f4",
X"a3",
X"02",
X"00",
X"78",
X"a6",
X"03",
X"c4",
X"9c",
X"02",
X"03",
X"23",
X"02",
X"25",
X"02",
X"26",
X"02",
X"24",
X"02",
X"27",
X"02",
X"1d",
X"02",
X"1f",
X"02",
X"1e",
X"02",
X"20",
X"02",
X"21",
X"02",
X"22",
X"02",
X"2a",
X"02",
X"29",
X"03",
X"01",
X"1f",
X"a3",
X"c2",
X"03",
X"0d",
X"2b",
X"0f",
X"38",
X"0e",
X"c4",
X"2c",
X"02",
X"03",
X"12",
X"0f",
X"3c",
X"0e",
X"02",
X"03",
X"44",
X"d2",
X"02",
X"00",
X"c8",
X"a7",
X"d3",
X"02",
X"c2",
X"03",
X"3f",
X"2b",
X"0f",
X"3a",
X"00",
X"d4",
X"a7",
X"2c",
X"03",
X"2b",
X"0f",
X"3a",
X"0e",
X"2c",
X"03",
X"2b",
X"0f",
X"3a",
X"c7",
X"2c",
X"03",
X"c4",
X"e3",
X"c2",
X"03",
X"c8",
X"02",
X"cb",
X"02",
X"01",
X"1b",
X"a4",
X"03",
X"00",
X"d0",
X"a7",
X"a5",
X"03",
X"01",
X"23",
X"a3",
X"c2",
X"03",
X"2b",
X"0f",
X"37",
X"0e",
X"c4",
X"2c",
X"02",
X"03",
X"12",
X"0f",
X"3c",
X"0e",
X"02",
X"03",
X"1d",
X"0f",
X"2f",
X"02",
X"1e",
X"0f",
X"30",
X"02",
X"1f",
X"0f",
X"31",
X"02",
X"20",
X"0f",
X"32",
X"02",
X"21",
X"0f",
X"33",
X"02",
X"22",
X"0f",
X"34",
X"03",
X"1c",
X"0e",
X"12",
X"0e",
X"fa",
X"03",
X"00",
X"45",
X"a6",
X"22",
X"0f",
X"2d",
X"0e",
X"f1",
X"02",
X"86",
X"22",
X"0f",
X"2e",
X"00",
X"7c",
X"a6",
X"e8",
X"03",
X"01",
X"1f",
X"a3",
X"22",
X"0f",
X"2d",
X"0e",
X"19",
X"0e",
X"c3",
X"dc",
X"03",
X"1a",
X"0e",
X"02",
X"03",
X"0e",
X"12",
X"0e",
X"12",
X"c4",
X"03",
X"dd",
X"12",
X"01",
X"1f",
X"a3",
X"cb",
X"03",
X"0e",
X"c8",
X"02",
X"c6",
X"03",
X"f7",
X"db",
X"c2",
X"03",
X"14",
X"02",
X"16",
X"03",
X"c9",
X"bb",
X"02",
X"ec",
X"00",
X"9a",
X"a7",
X"b5",
X"03",
X"1c",
X"0e",
X"03",
X"01",
X"1f",
X"a3",
X"02",
X"01",
X"23",
X"a3",
X"03",
X"b8",
X"c2",
X"03",
X"12",
X"bc",
X"02",
X"03",
X"0e",
X"12",
X"ac",
X"12",
X"f9",
X"12",
X"f3",
X"9a",
X"03",
X"a5",
X"97",
X"03",
X"ed",
X"94",
X"03",
X"ea",
X"91",
X"02",
X"8f",
X"03",
X"9a",
X"12",
X"02",
X"97",
X"15",
X"02",
X"03",
X"de",
X"85",
X"02",
X"db",
X"12",
X"c4",
X"02",
X"c2",
X"03",
X"00",
X"ba",
X"a7",
X"f4",
X"03",
X"c3",
X"f1",
X"03",
X"82",
X"12",
X"00",
X"45",
X"a6",
X"03",
X"ba",
X"12",
X"00",
X"45",
X"a6",
X"e4",
X"03",
X"00",
X"7c",
X"a6",
X"03",
X"0e",
X"12",
X"0e",
X"03",
X"0e",
X"12",
X"0e",
X"12",
X"b8",
X"d5",
X"03",
X"ed",
X"d2",
X"03",
X"0e",
X"c4",
X"c7",
X"cd",
X"03",
X"17",
X"02",
X"18",
X"03",
X"0e",
X"c2",
X"03",
X"12",
X"bc",
X"02",
X"03",
X"14",
X"02",
X"16",
X"03",
X"01",
X"1f",
X"a3",
X"0d",
X"2b",
X"0f",
X"39",
X"0e",
X"00",
X"53",
X"a6",
X"2c",
X"02",
X"01",
X"23",
X"a3",
X"2b",
X"0f",
X"3b",
X"0e",
X"2c",
X"03",
X"aa",
X"c3",
X"02",
X"03",
X"12",
X"bb",
X"02",
X"03",
X"0e",
X"1b",
X"c3",
X"9b",
X"03",
X"01",
X"f4",
X"a3",
X"02",
X"01",
X"ce",
X"a2",
X"c9",
X"02",
X"d4",
X"c3",
X"02",
X"03",
X"c3",
X"02",
X"03",
X"c3",
X"c8",
X"03",
X"0e",
X"02",
X"00",
X"7c",
X"a6",
X"03",
X"c4",
X"b3",
X"02",
X"03",
X"c6",
X"c2",
X"03",
X"bd",
X"02",
X"03",
X"12",
X"02",
X"15",
X"03",
X"0e",
X"c3",
X"02",
X"03",
X"12",
X"0e",
X"02",
X"03",
X"01",
X"da",
X"a2",
X"01",
X"da",
X"a2",
X"40",
X"02",
X"41",
X"02",
X"43",
X"02",
X"42",
X"03",
X"3d",
X"02",
X"3e",
X"03",
X"0e",
X"c2",
X"03",
X"12",
X"0f",
X"3c",
X"ba",
X"02",
X"03",
X"82",
X"80",
X"ac",
X"a4",
X"ba",
X"bb",
X"9b",
X"47",
X"4f",
X"54",
X"cf",
X"47",
X"4f",
X"53",
X"55",
X"c2",
X"54",
X"cf",
X"53",
X"54",
X"45",
X"d0",
X"54",
X"48",
X"45",
X"ce",
X"a3",
X"3c",
X"bd",
X"3c",
X"be",
X"3e",
X"bd",
X"bc",
X"be",
X"bd",
X"de",
X"aa",
X"ab",
X"ad",
X"af",
X"4e",
X"4f",
X"d4",
X"4f",
X"d2",
X"41",
X"4e",
X"c4",
X"a8",
X"a9",
X"bd",
X"bd",
X"3c",
X"bd",
X"3c",
X"be",
X"3e",
X"bd",
X"bc",
X"be",
X"bd",
X"ab",
X"ad",
X"a8",
X"80",
X"80",
X"a8",
X"a8",
X"ac",
X"53",
X"54",
X"52",
X"a4",
X"43",
X"48",
X"52",
X"a4",
X"55",
X"53",
X"d2",
X"41",
X"53",
X"c3",
X"56",
X"41",
X"cc",
X"4c",
X"45",
X"ce",
X"41",
X"44",
X"d2",
X"41",
X"54",
X"ce",
X"43",
X"4f",
X"d3",
X"50",
X"45",
X"45",
X"cb",
X"53",
X"49",
X"ce",
X"52",
X"4e",
X"c4",
X"46",
X"52",
X"c5",
X"45",
X"58",
X"d0",
X"4c",
X"4f",
X"c7",
X"43",
X"4c",
X"4f",
X"c7",
X"53",
X"51",
X"d2",
X"53",
X"47",
X"ce",
X"41",
X"42",
X"d3",
X"49",
X"4e",
X"d4",
X"50",
X"41",
X"44",
X"44",
X"4c",
X"c5",
X"53",
X"54",
X"49",
X"43",
X"cb",
X"50",
X"54",
X"52",
X"49",
X"c7",
X"53",
X"54",
X"52",
X"49",
X"c7",
X"00",
X"a9",
X"00",
X"84",
X"a4",
X"85",
X"a5",
X"98",
X"38",
X"65",
X"90",
X"a8",
X"a5",
X"91",
X"65",
X"a5",
X"cd",
X"e6",
X"02",
X"90",
X"0c",
X"d0",
X"07",
X"cc",
X"e5",
X"02",
X"90",
X"05",
X"f0",
X"03",
X"4c",
X"30",
X"b9",
X"38",
X"a5",
X"90",
X"f5",
X"00",
X"85",
X"a2",
X"a5",
X"91",
X"f5",
X"01",
X"85",
X"a3",
X"18",
X"75",
X"01",
X"85",
X"9a",
X"b5",
X"00",
X"85",
X"99",
X"85",
X"97",
X"65",
X"a4",
X"85",
X"9b",
X"b5",
X"01",
X"85",
X"98",
X"65",
X"a5",
X"65",
X"a3",
X"85",
X"9c",
X"b5",
X"00",
X"65",
X"a4",
X"95",
X"00",
X"b5",
X"01",
X"65",
X"a5",
X"95",
X"01",
X"e8",
X"e8",
X"e0",
X"92",
X"90",
X"ee",
X"85",
X"0f",
X"a5",
X"90",
X"85",
X"0e",
X"a6",
X"a3",
X"e8",
X"a4",
X"a2",
X"d0",
X"0d",
X"ea",
X"f0",
X"11",
X"ea",
X"88",
X"c6",
X"9a",
X"c6",
X"9c",
X"b1",
X"99",
X"91",
X"9b",
X"88",
X"d0",
X"f9",
X"b1",
X"99",
X"91",
X"9b",
X"ca",
X"d0",
X"ed",
X"60",
X"a8",
X"a9",
X"00",
X"84",
X"a4",
X"85",
X"a5",
X"38",
X"a5",
X"90",
X"f5",
X"00",
X"49",
X"ff",
X"a8",
X"c8",
X"84",
X"a2",
X"a5",
X"91",
X"f5",
X"01",
X"85",
X"a3",
X"b5",
X"00",
X"e5",
X"a2",
X"85",
X"99",
X"b5",
X"01",
X"e9",
X"00",
X"85",
X"9a",
X"86",
X"9b",
X"38",
X"b5",
X"00",
X"e5",
X"a4",
X"95",
X"00",
X"b5",
X"01",
X"e5",
X"a5",
X"95",
X"01",
X"e8",
X"e8",
X"e0",
X"92",
X"90",
X"ed",
X"85",
X"0f",
X"a5",
X"90",
X"85",
X"0e",
X"a6",
X"9b",
X"b5",
X"00",
X"e5",
X"a2",
X"85",
X"9b",
X"b5",
X"01",
X"e9",
X"00",
X"85",
X"9c",
X"a6",
X"a3",
X"e8",
X"a4",
X"a2",
X"d0",
X"08",
X"ca",
X"d0",
X"05",
X"60",
X"e6",
X"9a",
X"e6",
X"9c",
X"b1",
X"99",
X"91",
X"9b",
X"c8",
X"d0",
X"f9",
X"ca",
X"d0",
X"f2",
X"60",
X"20",
X"19",
X"b8",
X"20",
X"f2",
X"a9",
X"f0",
X"36",
X"a4",
X"a7",
X"c4",
X"9f",
X"b0",
X"1d",
X"b1",
X"8a",
X"85",
X"a7",
X"98",
X"c8",
X"b1",
X"8a",
X"c8",
X"84",
X"a8",
X"20",
X"7e",
X"a9",
X"ea",
X"4c",
X"61",
X"a9",
X"0a",
X"aa",
X"bd",
X"fa",
X"a9",
X"48",
X"bd",
X"fb",
X"a9",
X"48",
X"60",
X"a0",
X"01",
X"b1",
X"8a",
X"30",
X"10",
X"a5",
X"9f",
X"20",
X"d0",
X"a9",
X"20",
X"e1",
X"a9",
X"10",
X"c5",
X"4c",
X"8c",
X"b7",
X"4c",
X"92",
X"b7",
X"4c",
X"5d",
X"a0",
X"a5",
X"8a",
X"85",
X"be",
X"a5",
X"8b",
X"85",
X"bf",
X"a5",
X"89",
X"a4",
X"88",
X"85",
X"8b",
X"84",
X"8a",
X"a0",
X"01",
X"b1",
X"8a",
X"c5",
X"a1",
X"90",
X"0d",
X"d0",
X"0a",
X"88",
X"b1",
X"8a",
X"c5",
X"a0",
X"90",
X"04",
X"d0",
X"01",
X"18",
X"60",
X"20",
X"dc",
X"a9",
X"20",
X"d0",
X"a9",
X"4c",
X"b2",
X"a9",
X"18",
X"65",
X"8a",
X"85",
X"8a",
X"a5",
X"8b",
X"69",
X"00",
X"85",
X"8b",
X"60",
X"a0",
X"02",
X"b1",
X"8a",
X"60",
X"a0",
X"01",
X"b1",
X"8a",
X"60",
X"20",
X"45",
X"bd",
X"4c",
X"71",
X"e4",
X"20",
X"45",
X"bd",
X"6c",
X"0a",
X"00",
X"a4",
X"11",
X"d0",
X"03",
X"c6",
X"11",
X"98",
X"60",
X"a9",
X"e4",
X"a9",
X"e4",
X"b3",
X"3d",
X"ba",
X"1e",
X"b4",
X"b4",
X"ba",
X"c4",
X"aa",
X"d9",
X"b7",
X"77",
X"b6",
X"7c",
X"b6",
X"ff",
X"b6",
X"d4",
X"b6",
X"d4",
X"b6",
X"d1",
X"b7",
X"d7",
X"a9",
X"e5",
X"b7",
X"b4",
X"b2",
X"05",
X"bc",
X"21",
X"b7",
X"65",
X"b2",
X"8c",
X"b2",
X"05",
X"b7",
X"8b",
X"a0",
X"0b",
X"bb",
X"f1",
X"ba",
X"fa",
X"bb",
X"6c",
X"bc",
X"2e",
X"bc",
X"3c",
X"bc",
X"53",
X"bb",
X"eb",
X"b7",
X"e3",
X"b2",
X"77",
X"b3",
X"d9",
X"b2",
X"90",
X"b2",
X"ad",
X"b2",
X"95",
X"bd",
X"a7",
X"b7",
X"4b",
X"b7",
X"91",
X"b8",
X"3d",
X"b3",
X"d9",
X"bc",
X"84",
X"bc",
X"77",
X"ba",
X"45",
X"ba",
X"6b",
X"ba",
X"0b",
X"a9",
X"eb",
X"ba",
X"26",
X"b9",
X"ac",
X"bc",
X"9d",
X"b9",
X"d2",
X"b4",
X"95",
X"bb",
X"d0",
X"bb",
X"63",
X"aa",
X"d9",
X"b9",
X"11",
X"ac",
X"a2",
X"ac",
X"ab",
X"ac",
X"c1",
X"ac",
X"b1",
X"ac",
X"b8",
X"ac",
X"c8",
X"b1",
X"5d",
X"ac",
X"82",
X"bd",
X"f9",
X"ac",
X"79",
X"ac",
X"8b",
X"ac",
X"e3",
X"ac",
X"d8",
X"ac",
X"ce",
X"ab",
X"34",
X"ad",
X"65",
X"ad",
X"49",
X"ae",
X"8d",
X"ac",
X"a2",
X"ac",
X"ab",
X"ac",
X"c1",
X"ac",
X"b1",
X"ac",
X"b8",
X"ac",
X"c8",
X"ab",
X"34",
X"ac",
X"94",
X"ae",
X"10",
X"ad",
X"70",
X"ad",
X"6c",
X"ad",
X"65",
X"ad",
X"6c",
X"ad",
X"63",
X"b0",
X"33",
X"b0",
X"51",
X"b0",
X"a4",
X"af",
X"fc",
X"af",
X"ea",
X"af",
X"b4",
X"b0",
X"06",
X"b1",
X"17",
X"b1",
X"0e",
X"af",
X"cb",
X"b1",
X"05",
X"b0",
X"75",
X"af",
X"d5",
X"b1",
X"49",
X"b1",
X"20",
X"b1",
X"3c",
X"b1",
X"52",
X"ad",
X"03",
X"b0",
X"98",
X"b0",
X"c7",
X"b0",
X"0c",
X"b0",
X"10",
X"b0",
X"14",
X"b0",
X"18",
X"20",
X"26",
X"ab",
X"20",
X"36",
X"ab",
X"b0",
X"05",
X"20",
X"b2",
X"ab",
X"30",
X"f6",
X"85",
X"ab",
X"aa",
X"bd",
X"25",
X"ac",
X"4a",
X"4a",
X"4a",
X"4a",
X"85",
X"ac",
X"a4",
X"a9",
X"b1",
X"80",
X"aa",
X"bd",
X"25",
X"ac",
X"29",
X"0f",
X"c5",
X"ac",
X"90",
X"0d",
X"aa",
X"f0",
X"31",
X"b1",
X"80",
X"e6",
X"a9",
X"20",
X"18",
X"ab",
X"4c",
X"f3",
X"aa",
X"a5",
X"ab",
X"88",
X"91",
X"80",
X"84",
X"a9",
X"4c",
X"dd",
X"aa",
X"38",
X"e9",
X"1d",
X"0a",
X"aa",
X"bd",
X"6a",
X"aa",
X"48",
X"bd",
X"6b",
X"aa",
X"48",
X"60",
X"a0",
X"ff",
X"a9",
X"11",
X"91",
X"80",
X"84",
X"a9",
X"c8",
X"84",
X"b0",
X"84",
X"aa",
X"84",
X"b1",
X"60",
X"a4",
X"a8",
X"e6",
X"a8",
X"b1",
X"8a",
X"30",
X"43",
X"c9",
X"0f",
X"90",
X"03",
X"f0",
X"13",
X"60",
X"a2",
X"00",
X"c8",
X"b1",
X"8a",
X"95",
X"d4",
X"e8",
X"e0",
X"06",
X"90",
X"f6",
X"c8",
X"a9",
X"00",
X"aa",
X"f0",
X"22",
X"c8",
X"b1",
X"8a",
X"a2",
X"8a",
X"85",
X"d6",
X"85",
X"d8",
X"c8",
X"98",
X"18",
X"75",
X"00",
X"85",
X"d4",
X"a9",
X"00",
X"85",
X"d7",
X"85",
X"d9",
X"75",
X"01",
X"85",
X"d5",
X"98",
X"65",
X"d6",
X"a8",
X"a2",
X"00",
X"a9",
X"83",
X"85",
X"d2",
X"86",
X"d3",
X"84",
X"a8",
X"18",
X"60",
X"20",
X"1e",
X"ac",
X"b1",
X"9d",
X"99",
X"d2",
X"00",
X"c8",
X"c0",
X"08",
X"90",
X"f6",
X"18",
X"60",
X"20",
X"e9",
X"ab",
X"a9",
X"02",
X"24",
X"d2",
X"d0",
X"15",
X"05",
X"d2",
X"85",
X"d2",
X"6a",
X"90",
X"0f",
X"18",
X"a5",
X"d4",
X"65",
X"8c",
X"85",
X"d4",
X"a8",
X"a5",
X"d5",
X"65",
X"8d",
X"85",
X"d5",
X"60",
X"20",
X"22",
X"b9",
X"e6",
X"aa",
X"a5",
X"aa",
X"0a",
X"0a",
X"0a",
X"c5",
X"a9",
X"b0",
X"0d",
X"a8",
X"88",
X"a2",
X"07",
X"b5",
X"d2",
X"91",
X"80",
X"88",
X"ca",
X"10",
X"f8",
X"60",
X"4c",
X"20",
X"b9",
X"20",
X"d7",
X"ab",
X"a5",
X"d5",
X"10",
X"f5",
X"4c",
X"26",
X"b9",
X"20",
X"da",
X"aa",
X"20",
X"e9",
X"ab",
X"4c",
X"41",
X"ad",
X"20",
X"cd",
X"ab",
X"d0",
X"01",
X"60",
X"20",
X"2e",
X"b9",
X"a5",
X"aa",
X"c6",
X"aa",
X"0a",
X"0a",
X"0a",
X"a8",
X"88",
X"a2",
X"07",
X"b1",
X"80",
X"95",
X"d2",
X"88",
X"ca",
X"10",
X"f8",
X"60",
X"20",
X"e9",
X"ab",
X"20",
X"b6",
X"dd",
X"4c",
X"e9",
X"ab",
X"20",
X"da",
X"aa",
X"4c",
X"e9",
X"ab",
X"a5",
X"d3",
X"20",
X"1e",
X"ac",
X"a2",
X"00",
X"b5",
X"d2",
X"91",
X"9d",
X"c8",
X"e8",
X"e0",
X"08",
X"90",
X"f6",
X"60",
X"a0",
X"00",
X"84",
X"9e",
X"0a",
X"0a",
X"26",
X"9e",
X"0a",
X"26",
X"9e",
X"18",
X"65",
X"86",
X"85",
X"9d",
X"a5",
X"87",
X"65",
X"9e",
X"85",
X"9e",
X"60",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"88",
X"88",
X"88",
X"88",
X"88",
X"88",
X"cc",
X"aa",
X"99",
X"99",
X"aa",
X"dd",
X"55",
X"66",
X"f2",
X"4e",
X"f1",
X"f1",
X"ee",
X"ee",
X"ee",
X"ee",
X"ee",
X"ee",
X"dd",
X"dd",
X"f2",
X"f2",
X"f2",
X"f2",
X"f2",
X"43",
X"f2",
X"f2",
X"f2",
X"f2",
X"f2",
X"f2",
X"f2",
X"f2",
X"f2",
X"f2",
X"f2",
X"f2",
X"f2",
X"f2",
X"f2",
X"f2",
X"f2",
X"f2",
X"f2",
X"f2",
X"f2",
X"f2",
X"f2",
X"f2",
X"20",
X"fd",
X"ab",
X"20",
X"2c",
X"ad",
X"4c",
X"b2",
X"ab",
X"20",
X"fd",
X"ab",
X"20",
X"32",
X"ad",
X"4c",
X"b2",
X"ab",
X"20",
X"fd",
X"ab",
X"20",
X"38",
X"ad",
X"4c",
X"b2",
X"ab",
X"20",
X"e9",
X"ab",
X"a5",
X"d4",
X"f0",
X"04",
X"49",
X"80",
X"85",
X"d4",
X"4c",
X"b2",
X"ab",
X"20",
X"11",
X"ad",
X"30",
X"48",
X"f0",
X"46",
X"10",
X"3f",
X"20",
X"11",
X"ad",
X"4c",
X"e0",
X"ac",
X"20",
X"11",
X"ad",
X"30",
X"39",
X"10",
X"32",
X"20",
X"11",
X"ad",
X"30",
X"2d",
X"f0",
X"2b",
X"10",
X"2e",
X"20",
X"11",
X"ad",
X"30",
X"24",
X"10",
X"27",
X"20",
X"11",
X"ad",
X"4c",
X"e9",
X"ac",
X"20",
X"fd",
X"ab",
X"a5",
X"d4",
X"25",
X"e0",
X"4c",
X"e0",
X"ac",
X"20",
X"fd",
X"ab",
X"a5",
X"d4",
X"05",
X"e0",
X"f0",
X"09",
X"d0",
X"0c",
X"20",
X"e9",
X"ab",
X"a5",
X"d4",
X"f0",
X"05",
X"a9",
X"00",
X"a8",
X"f0",
X"04",
X"a9",
X"40",
X"a0",
X"01",
X"85",
X"d4",
X"84",
X"d5",
X"a2",
X"d6",
X"a0",
X"04",
X"20",
X"48",
X"da",
X"85",
X"d2",
X"4c",
X"b2",
X"ab",
X"20",
X"e9",
X"ab",
X"a5",
X"d4",
X"f0",
X"f6",
X"10",
X"e3",
X"a9",
X"c0",
X"30",
X"e1",
X"a4",
X"a9",
X"88",
X"b1",
X"80",
X"c9",
X"2f",
X"90",
X"03",
X"4c",
X"6c",
X"af",
X"20",
X"fd",
X"ab",
X"20",
X"2c",
X"ad",
X"a5",
X"d4",
X"60",
X"20",
X"66",
X"da",
X"b0",
X"13",
X"60",
X"20",
X"60",
X"da",
X"b0",
X"0d",
X"60",
X"20",
X"db",
X"da",
X"b0",
X"07",
X"60",
X"20",
X"28",
X"db",
X"b0",
X"01",
X"60",
X"20",
X"1e",
X"b9",
X"20",
X"d2",
X"d9",
X"b0",
X"01",
X"60",
X"20",
X"2e",
X"b9",
X"a5",
X"a9",
X"c9",
X"ff",
X"d0",
X"0f",
X"20",
X"fd",
X"ab",
X"a2",
X"05",
X"b5",
X"e0",
X"95",
X"d4",
X"ca",
X"10",
X"f9",
X"4c",
X"0c",
X"ac",
X"a9",
X"80",
X"85",
X"b1",
X"60",
X"e6",
X"b0",
X"a4",
X"a9",
X"68",
X"68",
X"4c",
X"04",
X"ab",
X"a9",
X"40",
X"85",
X"b1",
X"24",
X"b1",
X"10",
X"06",
X"a5",
X"aa",
X"85",
X"af",
X"c6",
X"aa",
X"a9",
X"00",
X"a8",
X"c5",
X"b0",
X"f0",
X"0b",
X"c6",
X"b0",
X"20",
X"da",
X"ab",
X"a5",
X"d5",
X"30",
X"23",
X"a4",
X"d4",
X"85",
X"98",
X"84",
X"97",
X"20",
X"da",
X"ab",
X"a5",
X"d4",
X"85",
X"f5",
X"a5",
X"d5",
X"30",
X"12",
X"85",
X"f6",
X"20",
X"e9",
X"ab",
X"24",
X"b1",
X"50",
X"05",
X"a9",
X"00",
X"85",
X"b1",
X"60",
X"66",
X"d2",
X"b0",
X"03",
X"20",
X"22",
X"b9",
X"a5",
X"f6",
X"c5",
X"d7",
X"90",
X"08",
X"d0",
X"f5",
X"a5",
X"f5",
X"c5",
X"d6",
X"b0",
X"ef",
X"a5",
X"98",
X"c5",
X"d9",
X"90",
X"08",
X"d0",
X"e7",
X"a5",
X"97",
X"c5",
X"d8",
X"b0",
X"e1",
X"20",
X"48",
X"af",
X"a5",
X"97",
X"a4",
X"98",
X"20",
X"3d",
X"af",
X"20",
X"31",
X"af",
X"a5",
X"d4",
X"a4",
X"d5",
X"20",
X"3d",
X"af",
X"a5",
X"8c",
X"a4",
X"8d",
X"20",
X"3d",
X"af",
X"24",
X"b1",
X"10",
X"15",
X"a5",
X"af",
X"85",
X"aa",
X"20",
X"e9",
X"ab",
X"a0",
X"05",
X"b9",
X"d4",
X"00",
X"91",
X"f5",
X"88",
X"10",
X"f8",
X"c8",
X"84",
X"b1",
X"60",
X"a0",
X"05",
X"b1",
X"f5",
X"99",
X"d4",
X"00",
X"88",
X"10",
X"f8",
X"c8",
X"84",
X"d2",
X"4c",
X"b2",
X"ab",
X"a5",
X"b0",
X"f0",
X"07",
X"20",
X"81",
X"ae",
X"84",
X"98",
X"85",
X"97",
X"20",
X"81",
X"ae",
X"38",
X"e9",
X"01",
X"85",
X"f5",
X"98",
X"e9",
X"00",
X"85",
X"f6",
X"20",
X"e9",
X"ab",
X"a5",
X"b1",
X"10",
X"0b",
X"05",
X"b0",
X"85",
X"b1",
X"a4",
X"d9",
X"a5",
X"d8",
X"4c",
X"3f",
X"ae",
X"a5",
X"d6",
X"a4",
X"d7",
X"a6",
X"b0",
X"f0",
X"10",
X"c6",
X"b0",
X"c4",
X"98",
X"90",
X"35",
X"d0",
X"04",
X"c5",
X"97",
X"90",
X"2f",
X"a4",
X"98",
X"a5",
X"97",
X"38",
X"e5",
X"f5",
X"85",
X"d6",
X"aa",
X"98",
X"e5",
X"f6",
X"85",
X"d7",
X"90",
X"1e",
X"a8",
X"d0",
X"03",
X"8a",
X"f0",
X"18",
X"20",
X"93",
X"ab",
X"18",
X"a5",
X"d4",
X"65",
X"f5",
X"85",
X"d4",
X"a5",
X"d5",
X"65",
X"f6",
X"85",
X"d5",
X"24",
X"b1",
X"10",
X"01",
X"60",
X"4c",
X"b2",
X"ab",
X"20",
X"2a",
X"b9",
X"20",
X"da",
X"ab",
X"a5",
X"d4",
X"a4",
X"d5",
X"d0",
X"03",
X"aa",
X"f0",
X"f1",
X"60",
X"20",
X"90",
X"ab",
X"a5",
X"d4",
X"85",
X"99",
X"a5",
X"d5",
X"85",
X"9a",
X"a5",
X"d6",
X"85",
X"a2",
X"a4",
X"d7",
X"84",
X"a3",
X"a4",
X"a9",
X"c0",
X"ff",
X"f0",
X"0f",
X"a9",
X"80",
X"85",
X"b1",
X"20",
X"04",
X"ab",
X"a5",
X"d7",
X"a4",
X"d6",
X"26",
X"b1",
X"b0",
X"07",
X"20",
X"90",
X"ab",
X"a5",
X"d9",
X"a4",
X"d8",
X"c5",
X"a3",
X"90",
X"06",
X"d0",
X"08",
X"c4",
X"a2",
X"b0",
X"04",
X"85",
X"a3",
X"84",
X"a2",
X"18",
X"a5",
X"d4",
X"65",
X"a2",
X"a8",
X"a5",
X"d5",
X"65",
X"a3",
X"aa",
X"38",
X"98",
X"e5",
X"8c",
X"85",
X"f9",
X"8a",
X"e5",
X"8d",
X"85",
X"fa",
X"38",
X"a9",
X"00",
X"e5",
X"a2",
X"85",
X"a2",
X"38",
X"a5",
X"99",
X"e5",
X"a2",
X"85",
X"99",
X"a5",
X"9a",
X"e9",
X"00",
X"85",
X"9a",
X"38",
X"a5",
X"d4",
X"e5",
X"a2",
X"85",
X"9b",
X"a5",
X"d5",
X"e9",
X"00",
X"85",
X"9c",
X"20",
X"44",
X"a9",
X"a5",
X"d3",
X"20",
X"81",
X"ab",
X"38",
X"a5",
X"f9",
X"e5",
X"d4",
X"a8",
X"a5",
X"fa",
X"e5",
X"d5",
X"aa",
X"a9",
X"02",
X"25",
X"b1",
X"f0",
X"0f",
X"a9",
X"00",
X"85",
X"b1",
X"e4",
X"d7",
X"90",
X"06",
X"d0",
X"05",
X"c4",
X"d6",
X"b0",
X"01",
X"60",
X"84",
X"d6",
X"86",
X"d7",
X"4c",
X"0c",
X"ac",
X"06",
X"f5",
X"26",
X"f6",
X"a4",
X"f6",
X"a5",
X"f5",
X"06",
X"f5",
X"26",
X"f6",
X"18",
X"65",
X"f5",
X"85",
X"f5",
X"98",
X"65",
X"f6",
X"85",
X"f6",
X"60",
X"a9",
X"00",
X"85",
X"f7",
X"85",
X"f8",
X"a0",
X"10",
X"a5",
X"f5",
X"4a",
X"90",
X"0c",
X"18",
X"a2",
X"fe",
X"b5",
X"f9",
X"75",
X"da",
X"95",
X"f9",
X"e8",
X"d0",
X"f7",
X"a2",
X"03",
X"76",
X"f5",
X"ca",
X"10",
X"fb",
X"88",
X"d0",
X"e5",
X"60",
X"20",
X"90",
X"ab",
X"20",
X"b6",
X"dd",
X"20",
X"90",
X"ab",
X"a2",
X"d6",
X"20",
X"a7",
X"af",
X"08",
X"a2",
X"e2",
X"20",
X"a7",
X"af",
X"f0",
X"13",
X"28",
X"f0",
X"0d",
X"a0",
X"00",
X"b1",
X"d4",
X"d1",
X"e0",
X"f0",
X"0c",
X"90",
X"03",
X"a9",
X"01",
X"60",
X"a9",
X"80",
X"60",
X"28",
X"d0",
X"f7",
X"60",
X"e6",
X"d4",
X"d0",
X"02",
X"e6",
X"d5",
X"e6",
X"e0",
X"d0",
X"d2",
X"e6",
X"e1",
X"d0",
X"ce",
X"b5",
X"00",
X"d0",
X"06",
X"b5",
X"01",
X"f0",
X"05",
X"d6",
X"01",
X"d6",
X"00",
X"a8",
X"60",
X"20",
X"90",
X"ab",
X"a5",
X"d6",
X"a4",
X"d7",
X"85",
X"d4",
X"84",
X"d5",
X"20",
X"aa",
X"d9",
X"a9",
X"00",
X"85",
X"d2",
X"85",
X"d3",
X"4c",
X"b2",
X"ab",
X"20",
X"da",
X"ab",
X"a0",
X"00",
X"b1",
X"d4",
X"4c",
X"bc",
X"af",
X"20",
X"e9",
X"ab",
X"38",
X"ad",
X"e5",
X"02",
X"e5",
X"90",
X"85",
X"d4",
X"ad",
X"e6",
X"02",
X"e5",
X"91",
X"85",
X"d5",
X"4c",
X"c0",
X"af",
X"20",
X"7d",
X"bd",
X"a9",
X"00",
X"85",
X"f2",
X"20",
X"00",
X"d8",
X"20",
X"9d",
X"bd",
X"90",
X"c9",
X"20",
X"10",
X"b9",
X"20",
X"90",
X"ab",
X"a0",
X"00",
X"b1",
X"d4",
X"4c",
X"bc",
X"af",
X"20",
X"90",
X"ab",
X"4c",
X"c0",
X"af",
X"a9",
X"00",
X"f0",
X"0a",
X"a9",
X"08",
X"d0",
X"06",
X"a9",
X"0c",
X"d0",
X"02",
X"a9",
X"14",
X"48",
X"20",
X"da",
X"ab",
X"a5",
X"d5",
X"d0",
X"0e",
X"a5",
X"d4",
X"68",
X"18",
X"65",
X"d4",
X"aa",
X"bd",
X"70",
X"02",
X"a0",
X"00",
X"f0",
X"8b",
X"20",
X"2e",
X"b9",
X"20",
X"e9",
X"ab",
X"20",
X"e6",
X"d8",
X"a5",
X"f3",
X"85",
X"d4",
X"a5",
X"f4",
X"85",
X"d5",
X"a0",
X"ff",
X"c8",
X"b1",
X"f3",
X"10",
X"fb",
X"29",
X"7f",
X"91",
X"f3",
X"c8",
X"84",
X"d6",
X"d0",
X"17",
X"20",
X"e9",
X"ab",
X"20",
X"41",
X"ad",
X"a5",
X"d4",
X"8d",
X"c0",
X"05",
X"a9",
X"05",
X"85",
X"d5",
X"a9",
X"c0",
X"85",
X"d4",
X"a9",
X"01",
X"85",
X"d6",
X"a9",
X"00",
X"85",
X"d7",
X"85",
X"d3",
X"a9",
X"83",
X"85",
X"d2",
X"4c",
X"b2",
X"ab",
X"a2",
X"93",
X"a0",
X"b0",
X"20",
X"98",
X"dd",
X"20",
X"e9",
X"ab",
X"ac",
X"0a",
X"d2",
X"84",
X"d4",
X"ac",
X"0a",
X"d2",
X"84",
X"d5",
X"20",
X"aa",
X"d9",
X"20",
X"38",
X"ad",
X"4c",
X"b2",
X"ab",
X"42",
X"06",
X"55",
X"36",
X"00",
X"00",
X"20",
X"e9",
X"ab",
X"a5",
X"d4",
X"29",
X"7f",
X"85",
X"d4",
X"4c",
X"b2",
X"ab",
X"20",
X"ae",
X"b0",
X"20",
X"aa",
X"d9",
X"4c",
X"b2",
X"ab",
X"a5",
X"b0",
X"85",
X"c6",
X"20",
X"da",
X"ab",
X"c6",
X"c6",
X"30",
X"09",
X"a5",
X"d4",
X"48",
X"a5",
X"d5",
X"48",
X"4c",
X"b2",
X"b0",
X"a5",
X"b0",
X"48",
X"6c",
X"d4",
X"00",
X"20",
X"e9",
X"ab",
X"20",
X"d1",
X"b0",
X"4c",
X"b2",
X"ab",
X"a5",
X"d4",
X"29",
X"7f",
X"38",
X"e9",
X"3f",
X"10",
X"02",
X"a9",
X"00",
X"aa",
X"a9",
X"00",
X"a8",
X"e0",
X"05",
X"b0",
X"07",
X"15",
X"d5",
X"94",
X"d5",
X"e8",
X"d0",
X"f5",
X"a6",
X"d4",
X"10",
X"14",
X"aa",
X"f0",
X"11",
X"a2",
X"e0",
X"20",
X"46",
X"da",
X"a9",
X"c0",
X"85",
X"e0",
X"a9",
X"01",
X"85",
X"e1",
X"20",
X"26",
X"ad",
X"60",
X"4c",
X"00",
X"dc",
X"20",
X"e9",
X"ab",
X"20",
X"05",
X"be",
X"4c",
X"59",
X"b1",
X"20",
X"e9",
X"ab",
X"20",
X"0f",
X"be",
X"4c",
X"59",
X"b1",
X"20",
X"e9",
X"ab",
X"20",
X"d5",
X"be",
X"4c",
X"59",
X"b1",
X"20",
X"e9",
X"ab",
X"a5",
X"d4",
X"f0",
X"33",
X"20",
X"cd",
X"de",
X"b0",
X"2e",
X"a5",
X"d4",
X"49",
X"3b",
X"d0",
X"39",
X"a5",
X"d5",
X"29",
X"f8",
X"d0",
X"33",
X"85",
X"d4",
X"f0",
X"2f",
X"20",
X"e9",
X"ab",
X"a5",
X"d4",
X"f0",
X"17",
X"20",
X"d1",
X"de",
X"4c",
X"2b",
X"b1",
X"20",
X"e9",
X"ab",
X"20",
X"c0",
X"dd",
X"4c",
X"59",
X"b1",
X"20",
X"e9",
X"ab",
X"20",
X"43",
X"bf",
X"90",
X"11",
X"20",
X"2e",
X"b9",
X"20",
X"fd",
X"ab",
X"a5",
X"e0",
X"f0",
X"0a",
X"2a",
X"a4",
X"d4",
X"d0",
X"08",
X"b0",
X"ef",
X"4c",
X"b2",
X"ab",
X"4c",
X"f0",
X"ac",
X"a2",
X"d4",
X"20",
X"76",
X"ba",
X"6a",
X"48",
X"a2",
X"e0",
X"20",
X"76",
X"ba",
X"98",
X"10",
X"1e",
X"29",
X"7f",
X"85",
X"d4",
X"b0",
X"03",
X"68",
X"90",
X"d1",
X"a5",
X"e0",
X"10",
X"01",
X"18",
X"08",
X"a6",
X"f7",
X"e0",
X"05",
X"b0",
X"0f",
X"b5",
X"e1",
X"6a",
X"90",
X"0a",
X"a9",
X"80",
X"d0",
X"08",
X"a5",
X"e0",
X"10",
X"01",
X"18",
X"08",
X"a9",
X"00",
X"48",
X"a2",
X"05",
X"b5",
X"e0",
X"48",
X"ca",
X"10",
X"fa",
X"20",
X"d1",
X"de",
X"a2",
X"00",
X"a0",
X"05",
X"68",
X"95",
X"e0",
X"e8",
X"88",
X"10",
X"f9",
X"20",
X"32",
X"ad",
X"20",
X"cc",
X"dd",
X"b0",
X"3d",
X"68",
X"05",
X"d4",
X"85",
X"d4",
X"28",
X"68",
X"10",
X"9d",
X"90",
X"9b",
X"a2",
X"d4",
X"20",
X"76",
X"ba",
X"b0",
X"94",
X"a5",
X"d4",
X"38",
X"29",
X"7f",
X"e9",
X"3f",
X"c9",
X"06",
X"b0",
X"1d",
X"aa",
X"a8",
X"f8",
X"38",
X"b5",
X"d4",
X"69",
X"00",
X"95",
X"d4",
X"ca",
X"d0",
X"f7",
X"d8",
X"90",
X"04",
X"e6",
X"d4",
X"e6",
X"d5",
X"c8",
X"c0",
X"06",
X"b0",
X"04",
X"96",
X"d4",
X"90",
X"f7",
X"4c",
X"b2",
X"ab",
X"20",
X"1e",
X"b9",
X"a4",
X"a8",
X"c4",
X"a7",
X"90",
X"01",
X"60",
X"20",
X"da",
X"aa",
X"a5",
X"d2",
X"6a",
X"90",
X"03",
X"20",
X"22",
X"b9",
X"38",
X"2a",
X"85",
X"d2",
X"30",
X"2e",
X"a4",
X"f5",
X"a6",
X"f6",
X"c8",
X"d0",
X"03",
X"e8",
X"30",
X"ed",
X"84",
X"d6",
X"86",
X"d7",
X"84",
X"f5",
X"86",
X"f6",
X"a4",
X"97",
X"a6",
X"98",
X"c8",
X"d0",
X"03",
X"e8",
X"30",
X"db",
X"84",
X"d8",
X"86",
X"d9",
X"20",
X"48",
X"af",
X"20",
X"31",
X"af",
X"a4",
X"f5",
X"a5",
X"f6",
X"30",
X"cb",
X"10",
X"14",
X"a9",
X"00",
X"85",
X"d6",
X"85",
X"d7",
X"a4",
X"f5",
X"84",
X"d8",
X"a5",
X"f6",
X"85",
X"d9",
X"d0",
X"04",
X"c0",
X"00",
X"f0",
X"b5",
X"a2",
X"8e",
X"20",
X"7c",
X"a8",
X"38",
X"a5",
X"97",
X"e5",
X"8c",
X"85",
X"d4",
X"a5",
X"98",
X"e5",
X"8d",
X"85",
X"d5",
X"20",
X"0c",
X"ac",
X"4c",
X"06",
X"b2",
X"20",
X"d7",
X"ab",
X"a5",
X"d4",
X"85",
X"95",
X"a5",
X"d5",
X"85",
X"96",
X"20",
X"e0",
X"ab",
X"a5",
X"d4",
X"a0",
X"00",
X"91",
X"95",
X"60",
X"a9",
X"06",
X"d0",
X"02",
X"a9",
X"00",
X"85",
X"fb",
X"60",
X"a9",
X"00",
X"85",
X"b6",
X"20",
X"04",
X"b9",
X"90",
X"03",
X"a8",
X"f0",
X"07",
X"20",
X"cd",
X"ab",
X"a5",
X"d5",
X"a4",
X"d4",
X"85",
X"b8",
X"84",
X"b7",
X"60",
X"a5",
X"a8",
X"48",
X"20",
X"f9",
X"b6",
X"a5",
X"b7",
X"85",
X"a0",
X"a5",
X"b8",
X"85",
X"a1",
X"20",
X"a2",
X"a9",
X"a5",
X"8a",
X"85",
X"f3",
X"a5",
X"8b",
X"85",
X"f4",
X"20",
X"a8",
X"bd",
X"68",
X"85",
X"a8",
X"a0",
X"00",
X"84",
X"f2",
X"20",
X"2f",
X"b3",
X"85",
X"b7",
X"20",
X"2d",
X"b3",
X"85",
X"b8",
X"20",
X"2d",
X"b3",
X"85",
X"f5",
X"20",
X"2d",
X"b3",
X"85",
X"f6",
X"20",
X"2d",
X"b3",
X"49",
X"01",
X"f0",
X"26",
X"a4",
X"f6",
X"c4",
X"f5",
X"b0",
X"05",
X"88",
X"84",
X"f2",
X"90",
X"e9",
X"84",
X"f2",
X"c6",
X"f2",
X"a0",
X"01",
X"b1",
X"f3",
X"30",
X"3a",
X"38",
X"a5",
X"f2",
X"65",
X"f3",
X"85",
X"f3",
X"a9",
X"00",
X"85",
X"b6",
X"65",
X"f4",
X"85",
X"f4",
X"90",
X"bb",
X"85",
X"f5",
X"a5",
X"f5",
X"c5",
X"b6",
X"b0",
X"0b",
X"20",
X"2d",
X"b3",
X"d0",
X"fb",
X"b0",
X"da",
X"e6",
X"f5",
X"d0",
X"ef",
X"a9",
X"40",
X"85",
X"a6",
X"e6",
X"f2",
X"b0",
X"32",
X"e6",
X"f2",
X"a4",
X"f2",
X"b1",
X"f3",
X"c9",
X"2c",
X"18",
X"f0",
X"02",
X"c9",
X"9b",
X"60",
X"20",
X"28",
X"b9",
X"a9",
X"3f",
X"85",
X"c2",
X"20",
X"36",
X"ab",
X"c6",
X"a8",
X"90",
X"05",
X"20",
X"07",
X"bd",
X"85",
X"b4",
X"20",
X"51",
X"da",
X"20",
X"e4",
X"bd",
X"20",
X"f2",
X"a9",
X"f0",
X"1f",
X"a0",
X"00",
X"84",
X"a6",
X"84",
X"f2",
X"20",
X"36",
X"ab",
X"e6",
X"a8",
X"a5",
X"d2",
X"30",
X"1a",
X"20",
X"00",
X"d8",
X"b0",
X"0e",
X"20",
X"2f",
X"b3",
X"d0",
X"09",
X"20",
X"0c",
X"ac",
X"4c",
X"ad",
X"b3",
X"4c",
X"92",
X"b7",
X"a9",
X"00",
X"85",
X"b4",
X"20",
X"24",
X"b9",
X"20",
X"26",
X"ab",
X"20",
X"b2",
X"ab",
X"c6",
X"f2",
X"a5",
X"f2",
X"85",
X"f5",
X"a2",
X"ff",
X"e8",
X"20",
X"2d",
X"b3",
X"d0",
X"fa",
X"b0",
X"04",
X"24",
X"a6",
X"50",
X"f4",
X"a4",
X"f5",
X"a5",
X"a8",
X"48",
X"8a",
X"a2",
X"f3",
X"20",
X"5c",
X"ab",
X"68",
X"85",
X"a8",
X"20",
X"91",
X"ae",
X"24",
X"a6",
X"50",
X"0f",
X"e6",
X"b6",
X"20",
X"04",
X"b9",
X"b0",
X"0d",
X"20",
X"2f",
X"b3",
X"90",
X"18",
X"4c",
X"fb",
X"b2",
X"20",
X"04",
X"b9",
X"90",
X"08",
X"20",
X"51",
X"da",
X"a9",
X"00",
X"85",
X"b4",
X"60",
X"20",
X"2f",
X"b3",
X"90",
X"03",
X"4c",
X"4e",
X"b3",
X"e6",
X"f2",
X"4c",
X"5f",
X"b3",
X"a5",
X"c9",
X"85",
X"af",
X"a9",
X"00",
X"85",
X"94",
X"a4",
X"a8",
X"b1",
X"8a",
X"c9",
X"12",
X"f0",
X"5f",
X"c9",
X"16",
X"f0",
X"79",
X"c9",
X"14",
X"f0",
X"75",
X"c9",
X"15",
X"f0",
X"7e",
X"c9",
X"1c",
X"f0",
X"70",
X"20",
X"da",
X"aa",
X"20",
X"e9",
X"ab",
X"c6",
X"a8",
X"24",
X"d2",
X"30",
X"22",
X"a5",
X"d5",
X"c9",
X"10",
X"90",
X"06",
X"a5",
X"d9",
X"29",
X"f0",
X"85",
X"d9",
X"20",
X"e6",
X"d8",
X"a9",
X"00",
X"85",
X"f2",
X"a4",
X"f2",
X"b1",
X"f3",
X"48",
X"e6",
X"f2",
X"20",
X"8f",
X"b4",
X"68",
X"10",
X"f3",
X"30",
X"ba",
X"20",
X"93",
X"ab",
X"a9",
X"00",
X"85",
X"f2",
X"a5",
X"d6",
X"d0",
X"04",
X"c6",
X"d7",
X"30",
X"ab",
X"c6",
X"d6",
X"a4",
X"f2",
X"b1",
X"d4",
X"e6",
X"f2",
X"d0",
X"02",
X"e6",
X"d5",
X"20",
X"91",
X"b4",
X"4c",
X"2f",
X"b4",
X"a4",
X"94",
X"c8",
X"c4",
X"af",
X"90",
X"09",
X"18",
X"a5",
X"c9",
X"65",
X"af",
X"85",
X"af",
X"90",
X"f0",
X"a4",
X"94",
X"c4",
X"af",
X"b0",
X"15",
X"a9",
X"20",
X"20",
X"8f",
X"b4",
X"4c",
X"59",
X"b4",
X"4c",
X"85",
X"b4",
X"20",
X"07",
X"bd",
X"85",
X"b5",
X"c6",
X"a8",
X"4c",
X"e2",
X"b3",
X"e6",
X"a8",
X"a4",
X"a8",
X"b1",
X"8a",
X"c9",
X"16",
X"f0",
X"0c",
X"c9",
X"14",
X"f0",
X"08",
X"4c",
X"e2",
X"b3",
X"a9",
X"9b",
X"20",
X"91",
X"b4",
X"a9",
X"00",
X"85",
X"b5",
X"60",
X"29",
X"7f",
X"e6",
X"94",
X"4c",
X"99",
X"ba",
X"a9",
X"b2",
X"85",
X"f3",
X"a9",
X"b4",
X"85",
X"f4",
X"a2",
X"07",
X"86",
X"b5",
X"a9",
X"00",
X"a0",
X"08",
X"20",
X"d8",
X"bb",
X"20",
X"bb",
X"bc",
X"20",
X"da",
X"b3",
X"4c",
X"f7",
X"bc",
X"50",
X"3a",
X"9b",
X"a0",
X"00",
X"84",
X"a0",
X"84",
X"a1",
X"88",
X"84",
X"ad",
X"a9",
X"7f",
X"85",
X"ae",
X"8d",
X"fe",
X"02",
X"a9",
X"9b",
X"20",
X"99",
X"ba",
X"20",
X"f9",
X"b6",
X"a4",
X"a8",
X"c8",
X"c4",
X"a7",
X"b0",
X"2d",
X"a5",
X"a8",
X"48",
X"20",
X"06",
X"ac",
X"68",
X"85",
X"a8",
X"a5",
X"d2",
X"10",
X"06",
X"20",
X"cf",
X"ba",
X"4c",
X"cd",
X"b4",
X"20",
X"cd",
X"ab",
X"85",
X"a1",
X"a5",
X"d4",
X"85",
X"a0",
X"a4",
X"a8",
X"c4",
X"a7",
X"f0",
X"03",
X"20",
X"cd",
X"ab",
X"a5",
X"d4",
X"85",
X"ad",
X"a5",
X"d5",
X"85",
X"ae",
X"20",
X"a2",
X"a9",
X"20",
X"e1",
X"a9",
X"30",
X"24",
X"a0",
X"01",
X"b1",
X"8a",
X"c5",
X"ae",
X"90",
X"0b",
X"d0",
X"1a",
X"88",
X"b1",
X"8a",
X"c5",
X"ad",
X"90",
X"02",
X"d0",
X"11",
X"20",
X"8e",
X"b5",
X"20",
X"f2",
X"a9",
X"f0",
X"09",
X"20",
X"dc",
X"a9",
X"20",
X"d0",
X"a9",
X"4c",
X"04",
X"b5",
X"a5",
X"b5",
X"f0",
X"07",
X"20",
X"f7",
X"bc",
X"a9",
X"00",
X"85",
X"b5",
X"8d",
X"fe",
X"02",
X"4c",
X"a8",
X"bd",
X"86",
X"aa",
X"20",
X"62",
X"b5",
X"a4",
X"aa",
X"c6",
X"af",
X"30",
X"0e",
X"b1",
X"95",
X"30",
X"03",
X"c8",
X"d0",
X"f9",
X"c8",
X"20",
X"57",
X"b5",
X"4c",
X"43",
X"b5",
X"18",
X"98",
X"65",
X"95",
X"85",
X"95",
X"a8",
X"a5",
X"96",
X"69",
X"00",
X"85",
X"96",
X"84",
X"95",
X"60",
X"a0",
X"ff",
X"84",
X"af",
X"e6",
X"af",
X"a4",
X"af",
X"b1",
X"95",
X"48",
X"c9",
X"9b",
X"f0",
X"04",
X"29",
X"7f",
X"f0",
X"03",
X"20",
X"99",
X"ba",
X"68",
X"10",
X"eb",
X"60",
X"a9",
X"20",
X"20",
X"99",
X"ba",
X"20",
X"67",
X"b5",
X"a9",
X"20",
X"4c",
X"99",
X"ba",
X"a0",
X"00",
X"b1",
X"8a",
X"85",
X"d4",
X"c8",
X"b1",
X"8a",
X"85",
X"d5",
X"20",
X"aa",
X"d9",
X"20",
X"e6",
X"d8",
X"a5",
X"f3",
X"85",
X"95",
X"a5",
X"f4",
X"85",
X"96",
X"20",
X"86",
X"b5",
X"a0",
X"02",
X"b1",
X"8a",
X"85",
X"9f",
X"c8",
X"b1",
X"8a",
X"85",
X"a7",
X"c8",
X"84",
X"a8",
X"20",
X"c2",
X"b5",
X"a4",
X"a7",
X"c4",
X"9f",
X"90",
X"f0",
X"60",
X"20",
X"63",
X"b6",
X"c9",
X"36",
X"f0",
X"17",
X"20",
X"6f",
X"b6",
X"20",
X"63",
X"b6",
X"c9",
X"37",
X"f0",
X"04",
X"c9",
X"02",
X"b0",
X"09",
X"20",
X"61",
X"b6",
X"20",
X"99",
X"ba",
X"4c",
X"d7",
X"b5",
X"20",
X"61",
X"b6",
X"10",
X"1a",
X"29",
X"7f",
X"85",
X"af",
X"a2",
X"00",
X"a5",
X"83",
X"a4",
X"82",
X"20",
X"3e",
X"b5",
X"20",
X"67",
X"b5",
X"c9",
X"a8",
X"d0",
X"e7",
X"20",
X"61",
X"b6",
X"4c",
X"e0",
X"b5",
X"c9",
X"0f",
X"f0",
X"18",
X"b0",
X"36",
X"20",
X"45",
X"ab",
X"c6",
X"a8",
X"20",
X"e6",
X"d8",
X"a5",
X"f3",
X"85",
X"95",
X"a5",
X"f4",
X"85",
X"96",
X"20",
X"67",
X"b5",
X"4c",
X"e0",
X"b5",
X"20",
X"61",
X"b6",
X"85",
X"af",
X"a9",
X"22",
X"20",
X"99",
X"ba",
X"a5",
X"af",
X"f0",
X"0a",
X"20",
X"61",
X"b6",
X"20",
X"99",
X"ba",
X"c6",
X"af",
X"d0",
X"f6",
X"a9",
X"22",
X"20",
X"99",
X"ba",
X"4c",
X"e0",
X"b5",
X"38",
X"e9",
X"10",
X"85",
X"af",
X"a2",
X"00",
X"a9",
X"a7",
X"a0",
X"de",
X"20",
X"3e",
X"b5",
X"20",
X"63",
X"b6",
X"c9",
X"3d",
X"b0",
X"c5",
X"a0",
X"00",
X"b1",
X"95",
X"29",
X"7f",
X"20",
X"ec",
X"a3",
X"b0",
X"ba",
X"20",
X"81",
X"b5",
X"4c",
X"e0",
X"b5",
X"e6",
X"a8",
X"a4",
X"a8",
X"c4",
X"a7",
X"b0",
X"03",
X"b1",
X"8a",
X"60",
X"68",
X"68",
X"60",
X"85",
X"af",
X"a2",
X"02",
X"a9",
X"a4",
X"a0",
X"9f",
X"20",
X"3e",
X"b5",
X"4c",
X"86",
X"b5",
X"20",
X"83",
X"b8",
X"20",
X"da",
X"aa",
X"a5",
X"d3",
X"09",
X"80",
X"48",
X"20",
X"23",
X"b8",
X"a9",
X"0c",
X"20",
X"71",
X"b8",
X"20",
X"06",
X"ac",
X"a2",
X"d4",
X"a0",
X"00",
X"20",
X"88",
X"b8",
X"20",
X"44",
X"da",
X"a9",
X"01",
X"85",
X"d5",
X"a9",
X"40",
X"85",
X"d4",
X"20",
X"04",
X"b9",
X"b0",
X"03",
X"20",
X"06",
X"ac",
X"a2",
X"d4",
X"a0",
X"06",
X"20",
X"88",
X"b8",
X"68",
X"48",
X"a9",
X"04",
X"20",
X"71",
X"b8",
X"68",
X"a0",
X"00",
X"91",
X"c4",
X"b1",
X"8a",
X"c8",
X"91",
X"c4",
X"b1",
X"8a",
X"c8",
X"91",
X"c4",
X"a6",
X"b3",
X"ca",
X"8a",
X"c8",
X"91",
X"c4",
X"60",
X"20",
X"f9",
X"b6",
X"20",
X"cd",
X"ab",
X"a5",
X"d5",
X"85",
X"a1",
X"a5",
X"d4",
X"85",
X"a0",
X"20",
X"a2",
X"a9",
X"b0",
X"05",
X"68",
X"68",
X"4c",
X"5e",
X"a9",
X"20",
X"f0",
X"b6",
X"20",
X"1c",
X"b9",
X"a5",
X"be",
X"85",
X"8a",
X"a5",
X"bf",
X"85",
X"8b",
X"60",
X"20",
X"83",
X"b8",
X"a9",
X"00",
X"f0",
X"b5",
X"a4",
X"a8",
X"b1",
X"8a",
X"85",
X"c7",
X"20",
X"3e",
X"b8",
X"b0",
X"3e",
X"f0",
X"3c",
X"c5",
X"c7",
X"d0",
X"f5",
X"a0",
X"06",
X"20",
X"97",
X"b8",
X"a5",
X"e0",
X"48",
X"a5",
X"c7",
X"20",
X"81",
X"ab",
X"20",
X"26",
X"ad",
X"20",
X"0c",
X"ac",
X"a0",
X"00",
X"20",
X"97",
X"b8",
X"68",
X"10",
X"06",
X"20",
X"20",
X"ad",
X"10",
X"09",
X"60",
X"20",
X"20",
X"ad",
X"f0",
X"03",
X"30",
X"01",
X"60",
X"a9",
X"10",
X"20",
X"71",
X"b8",
X"20",
X"cb",
X"bd",
X"c9",
X"08",
X"f0",
X"f3",
X"4c",
X"c2",
X"bd",
X"20",
X"1a",
X"b9",
X"20",
X"04",
X"b9",
X"b0",
X"03",
X"20",
X"f7",
X"ba",
X"ea",
X"a9",
X"00",
X"85",
X"a0",
X"85",
X"a1",
X"20",
X"16",
X"b8",
X"20",
X"e1",
X"a9",
X"30",
X"12",
X"20",
X"f1",
X"b8",
X"20",
X"b9",
X"b8",
X"20",
X"a8",
X"b8",
X"a9",
X"00",
X"85",
X"b7",
X"85",
X"b8",
X"85",
X"b6",
X"60",
X"4c",
X"50",
X"a0",
X"20",
X"06",
X"ac",
X"a5",
X"d5",
X"f0",
X"08",
X"20",
X"04",
X"b9",
X"b0",
X"07",
X"4c",
X"d5",
X"b6",
X"a5",
X"9f",
X"85",
X"a7",
X"60",
X"20",
X"a6",
X"b7",
X"4c",
X"50",
X"a0",
X"20",
X"a6",
X"b7",
X"20",
X"79",
X"bd",
X"a9",
X"fd",
X"85",
X"95",
X"a9",
X"a5",
X"85",
X"96",
X"20",
X"67",
X"b5",
X"4c",
X"68",
X"b9",
X"20",
X"e1",
X"a9",
X"30",
X"07",
X"85",
X"bb",
X"88",
X"b1",
X"8a",
X"85",
X"ba",
X"4c",
X"5b",
X"bd",
X"20",
X"e1",
X"a9",
X"10",
X"f8",
X"a5",
X"ba",
X"85",
X"a0",
X"a5",
X"bb",
X"85",
X"a1",
X"20",
X"a2",
X"a9",
X"20",
X"e1",
X"a9",
X"30",
X"ab",
X"20",
X"dc",
X"a9",
X"20",
X"d0",
X"a9",
X"20",
X"e1",
X"a9",
X"30",
X"a0",
X"4c",
X"19",
X"b8",
X"20",
X"d7",
X"ab",
X"a5",
X"d4",
X"85",
X"bc",
X"a5",
X"d5",
X"85",
X"bd",
X"60",
X"20",
X"83",
X"b8",
X"20",
X"e0",
X"ab",
X"a5",
X"d4",
X"f0",
X"23",
X"a4",
X"a8",
X"88",
X"b1",
X"8a",
X"c9",
X"17",
X"08",
X"f0",
X"03",
X"20",
X"fc",
X"b6",
X"a5",
X"d4",
X"85",
X"b3",
X"20",
X"cd",
X"ab",
X"c6",
X"b3",
X"f0",
X"0c",
X"20",
X"04",
X"b9",
X"90",
X"f4",
X"28",
X"f0",
X"03",
X"20",
X"3e",
X"b8",
X"60",
X"28",
X"4c",
X"d8",
X"b6",
X"20",
X"a2",
X"a9",
X"a0",
X"02",
X"b1",
X"8a",
X"85",
X"9f",
X"c8",
X"84",
X"a7",
X"60",
X"85",
X"c7",
X"20",
X"7a",
X"b8",
X"20",
X"3e",
X"b8",
X"b0",
X"08",
X"f0",
X"06",
X"c5",
X"c7",
X"f0",
X"0a",
X"d0",
X"f3",
X"a5",
X"c4",
X"85",
X"90",
X"a5",
X"c5",
X"85",
X"91",
X"60",
X"a5",
X"8f",
X"c5",
X"91",
X"90",
X"06",
X"a5",
X"8e",
X"c5",
X"90",
X"b0",
X"f3",
X"a9",
X"04",
X"a2",
X"90",
X"20",
X"f7",
X"a8",
X"a0",
X"03",
X"b1",
X"90",
X"85",
X"b2",
X"88",
X"b1",
X"90",
X"85",
X"a1",
X"88",
X"b1",
X"90",
X"85",
X"a0",
X"88",
X"b1",
X"90",
X"f0",
X"09",
X"48",
X"a9",
X"0c",
X"a2",
X"90",
X"20",
X"f7",
X"a8",
X"68",
X"18",
X"60",
X"20",
X"7a",
X"b8",
X"a8",
X"a2",
X"90",
X"4c",
X"7a",
X"a8",
X"a6",
X"90",
X"86",
X"c4",
X"a6",
X"91",
X"86",
X"c5",
X"60",
X"a4",
X"a8",
X"84",
X"b3",
X"60",
X"a9",
X"06",
X"85",
X"c6",
X"b5",
X"00",
X"91",
X"c4",
X"e8",
X"c8",
X"c6",
X"c6",
X"d0",
X"f6",
X"60",
X"a9",
X"06",
X"85",
X"c6",
X"a2",
X"e0",
X"b1",
X"90",
X"95",
X"00",
X"e8",
X"c8",
X"c6",
X"c6",
X"d0",
X"f6",
X"60",
X"a5",
X"8c",
X"85",
X"8e",
X"85",
X"90",
X"85",
X"0e",
X"a5",
X"8d",
X"85",
X"8f",
X"85",
X"91",
X"85",
X"0f",
X"60",
X"a6",
X"86",
X"86",
X"f5",
X"a4",
X"87",
X"84",
X"f6",
X"a6",
X"f6",
X"e4",
X"89",
X"90",
X"07",
X"a6",
X"f5",
X"e4",
X"88",
X"90",
X"01",
X"60",
X"a0",
X"00",
X"b1",
X"f5",
X"29",
X"fe",
X"91",
X"f5",
X"a0",
X"02",
X"a2",
X"06",
X"a9",
X"00",
X"91",
X"f5",
X"c8",
X"ca",
X"d0",
X"fa",
X"a5",
X"f5",
X"18",
X"69",
X"08",
X"85",
X"f5",
X"a5",
X"f6",
X"69",
X"00",
X"85",
X"f6",
X"d0",
X"d0",
X"a2",
X"05",
X"a0",
X"00",
X"94",
X"b6",
X"ca",
X"10",
X"fb",
X"84",
X"fb",
X"88",
X"84",
X"bd",
X"84",
X"11",
X"4c",
X"45",
X"bd",
X"a6",
X"a8",
X"e8",
X"e4",
X"a7",
X"60",
X"e6",
X"b9",
X"e6",
X"b9",
X"e6",
X"b9",
X"e6",
X"b9",
X"e6",
X"b9",
X"e6",
X"b9",
X"e6",
X"b9",
X"e6",
X"b9",
X"e6",
X"b9",
X"e6",
X"b9",
X"e6",
X"b9",
X"e6",
X"b9",
X"e6",
X"b9",
X"e6",
X"b9",
X"e6",
X"b9",
X"e6",
X"b9",
X"e6",
X"b9",
X"e6",
X"b9",
X"e6",
X"b9",
X"e6",
X"b9",
X"e6",
X"b9",
X"a9",
X"00",
X"8d",
X"fe",
X"02",
X"20",
X"a6",
X"b7",
X"a5",
X"bd",
X"30",
X"15",
X"85",
X"a1",
X"a5",
X"bc",
X"85",
X"a0",
X"a9",
X"80",
X"85",
X"bd",
X"a5",
X"b9",
X"85",
X"c3",
X"a9",
X"00",
X"85",
X"b9",
X"4c",
X"e0",
X"b6",
X"20",
X"79",
X"bd",
X"a9",
X"37",
X"20",
X"6f",
X"b6",
X"a5",
X"b9",
X"85",
X"d4",
X"a9",
X"00",
X"85",
X"d5",
X"20",
X"93",
X"b9",
X"20",
X"e1",
X"a9",
X"30",
X"19",
X"a9",
X"a4",
X"85",
X"95",
X"a9",
X"b9",
X"85",
X"96",
X"20",
X"67",
X"b5",
X"a0",
X"01",
X"b1",
X"8a",
X"85",
X"d5",
X"88",
X"b1",
X"8a",
X"85",
X"d4",
X"20",
X"93",
X"b9",
X"20",
X"79",
X"bd",
X"a9",
X"00",
X"85",
X"b9",
X"20",
X"5b",
X"bd",
X"4c",
X"60",
X"a0",
X"20",
X"aa",
X"d9",
X"20",
X"e6",
X"d8",
X"a5",
X"f3",
X"85",
X"95",
X"a5",
X"f4",
X"85",
X"96",
X"4c",
X"67",
X"b5",
X"20",
X"41",
X"54",
X"20",
X"4c",
X"49",
X"4e",
X"45",
X"a0",
X"20",
X"e0",
X"ab",
X"a5",
X"d4",
X"c9",
X"05",
X"b0",
X"1a",
X"48",
X"20",
X"d7",
X"ab",
X"a5",
X"d4",
X"0a",
X"0a",
X"0a",
X"0a",
X"48",
X"20",
X"d7",
X"ab",
X"68",
X"18",
X"65",
X"d4",
X"a8",
X"68",
X"aa",
X"98",
X"9d",
X"c4",
X"02",
X"60",
X"20",
X"2e",
X"b9",
X"20",
X"e0",
X"ab",
X"a5",
X"d4",
X"c9",
X"04",
X"b0",
X"f4",
X"0a",
X"48",
X"a9",
X"00",
X"8d",
X"08",
X"d2",
X"a9",
X"03",
X"8d",
X"0f",
X"d2",
X"20",
X"d7",
X"ab",
X"68",
X"48",
X"aa",
X"a5",
X"d4",
X"9d",
X"00",
X"d2",
X"20",
X"d7",
X"ab",
X"a5",
X"d4",
X"0a",
X"0a",
X"0a",
X"0a",
X"48",
X"20",
X"d7",
X"ab",
X"68",
X"a8",
X"68",
X"aa",
X"98",
X"18",
X"65",
X"d4",
X"9d",
X"01",
X"d2",
X"60",
X"20",
X"d7",
X"ab",
X"a5",
X"d4",
X"85",
X"55",
X"a5",
X"d5",
X"85",
X"56",
X"20",
X"e0",
X"ab",
X"a5",
X"d4",
X"85",
X"54",
X"60",
X"20",
X"d7",
X"ab",
X"a5",
X"d4",
X"85",
X"c8",
X"60",
X"20",
X"0c",
X"ba",
X"a5",
X"c8",
X"8d",
X"fb",
X"02",
X"a9",
X"11",
X"a2",
X"06",
X"20",
X"be",
X"ba",
X"a9",
X"0c",
X"9d",
X"4a",
X"03",
X"a9",
X"00",
X"9d",
X"4b",
X"03",
X"20",
X"29",
X"bd",
X"4c",
X"bb",
X"bc",
X"a2",
X"06",
X"86",
X"c1",
X"20",
X"f7",
X"bc",
X"20",
X"d7",
X"ab",
X"a2",
X"69",
X"a0",
X"ba",
X"86",
X"f3",
X"84",
X"f4",
X"a2",
X"06",
X"a5",
X"d4",
X"29",
X"f0",
X"49",
X"1c",
X"a8",
X"a5",
X"d4",
X"20",
X"d8",
X"bb",
X"4c",
X"bb",
X"bc",
X"53",
X"3a",
X"9b",
X"20",
X"0c",
X"ba",
X"a5",
X"c8",
X"a2",
X"06",
X"4c",
X"9b",
X"ba",
X"38",
X"b5",
X"00",
X"29",
X"7f",
X"e9",
X"40",
X"90",
X"19",
X"85",
X"f5",
X"85",
X"f7",
X"8a",
X"65",
X"f5",
X"e8",
X"e8",
X"e8",
X"e8",
X"e8",
X"e8",
X"86",
X"f5",
X"aa",
X"e8",
X"e4",
X"f5",
X"b0",
X"04",
X"b5",
X"00",
X"f0",
X"f7",
X"60",
X"a6",
X"b5",
X"48",
X"20",
X"c0",
X"ba",
X"bd",
X"4a",
X"03",
X"85",
X"2a",
X"bd",
X"4b",
X"03",
X"85",
X"2b",
X"68",
X"a8",
X"20",
X"b2",
X"ba",
X"98",
X"4c",
X"be",
X"bc",
X"bd",
X"47",
X"03",
X"48",
X"bd",
X"46",
X"03",
X"48",
X"98",
X"a0",
X"92",
X"60",
X"85",
X"c0",
X"86",
X"c1",
X"4c",
X"af",
X"bc",
X"a9",
X"04",
X"20",
X"d7",
X"ba",
X"85",
X"b4",
X"4c",
X"60",
X"a0",
X"a9",
X"08",
X"20",
X"d7",
X"ba",
X"85",
X"b5",
X"60",
X"48",
X"a0",
X"07",
X"84",
X"c1",
X"20",
X"af",
X"bc",
X"a9",
X"0c",
X"20",
X"2b",
X"bd",
X"a0",
X"03",
X"84",
X"c0",
X"68",
X"a0",
X"00",
X"20",
X"02",
X"bc",
X"a9",
X"07",
X"60",
X"40",
X"02",
X"00",
X"00",
X"00",
X"00",
X"a9",
X"ff",
X"d0",
X"02",
X"a9",
X"00",
X"48",
X"a9",
X"04",
X"20",
X"d7",
X"ba",
X"68",
X"48",
X"a9",
X"07",
X"85",
X"c0",
X"85",
X"ca",
X"20",
X"af",
X"bc",
X"a0",
X"0e",
X"20",
X"15",
X"bd",
X"20",
X"bb",
X"bc",
X"ad",
X"80",
X"05",
X"0d",
X"81",
X"05",
X"d0",
X"3f",
X"a2",
X"8c",
X"18",
X"a5",
X"80",
X"7d",
X"00",
X"05",
X"08",
X"18",
X"69",
X"00",
X"a8",
X"a5",
X"81",
X"7d",
X"01",
X"05",
X"28",
X"69",
X"00",
X"cd",
X"e6",
X"02",
X"90",
X"0a",
X"d0",
X"05",
X"cc",
X"e5",
X"02",
X"90",
X"03",
X"4c",
X"0e",
X"b9",
X"95",
X"01",
X"94",
X"00",
X"ca",
X"ca",
X"e0",
X"82",
X"b0",
X"d4",
X"20",
X"98",
X"bb",
X"20",
X"66",
X"b7",
X"a9",
X"00",
X"85",
X"ca",
X"68",
X"f0",
X"01",
X"60",
X"4c",
X"50",
X"a0",
X"a9",
X"00",
X"85",
X"ca",
X"20",
X"0a",
X"b9",
X"a9",
X"04",
X"20",
X"b4",
X"bb",
X"a9",
X"00",
X"f0",
X"97",
X"a9",
X"08",
X"20",
X"d7",
X"ba",
X"a9",
X"0b",
X"85",
X"c0",
X"a2",
X"80",
X"38",
X"b5",
X"00",
X"e5",
X"80",
X"9d",
X"00",
X"05",
X"e8",
X"b5",
X"00",
X"e5",
X"81",
X"9d",
X"00",
X"05",
X"e8",
X"e0",
X"8e",
X"90",
X"eb",
X"20",
X"af",
X"bc",
X"a0",
X"0e",
X"20",
X"15",
X"bd",
X"20",
X"bb",
X"bc",
X"20",
X"af",
X"bc",
X"a5",
X"82",
X"85",
X"f3",
X"a5",
X"83",
X"85",
X"f4",
X"ac",
X"8d",
X"05",
X"88",
X"98",
X"ac",
X"8c",
X"05",
X"20",
X"17",
X"bd",
X"20",
X"bb",
X"bc",
X"4c",
X"f7",
X"bc",
X"ea",
X"ea",
X"48",
X"a2",
X"ce",
X"86",
X"f3",
X"a2",
X"bb",
X"86",
X"f4",
X"a2",
X"07",
X"68",
X"a8",
X"a9",
X"80",
X"20",
X"d8",
X"bb",
X"20",
X"bb",
X"bc",
X"a9",
X"07",
X"60",
X"43",
X"3a",
X"9b",
X"a9",
X"08",
X"20",
X"b4",
X"bb",
X"d0",
X"9a",
X"48",
X"a9",
X"03",
X"20",
X"be",
X"ba",
X"68",
X"9d",
X"4b",
X"03",
X"98",
X"9d",
X"4a",
X"03",
X"20",
X"1e",
X"bd",
X"4c",
X"51",
X"da",
X"20",
X"09",
X"bd",
X"4c",
X"f4",
X"bb",
X"a9",
X"03",
X"85",
X"c0",
X"20",
X"a8",
X"bc",
X"20",
X"09",
X"bd",
X"48",
X"20",
X"09",
X"bd",
X"a8",
X"68",
X"48",
X"98",
X"48",
X"20",
X"da",
X"aa",
X"20",
X"7d",
X"bd",
X"20",
X"af",
X"bc",
X"68",
X"9d",
X"4b",
X"03",
X"68",
X"9d",
X"4a",
X"03",
X"20",
X"0f",
X"bd",
X"20",
X"9d",
X"bd",
X"20",
X"51",
X"da",
X"4c",
X"bb",
X"bc",
X"a9",
X"0c",
X"85",
X"c0",
X"20",
X"a8",
X"bc",
X"20",
X"29",
X"bd",
X"4c",
X"bb",
X"bc",
X"20",
X"a8",
X"bc",
X"a9",
X"0d",
X"20",
X"2b",
X"bd",
X"20",
X"00",
X"bd",
X"4c",
X"31",
X"bd",
X"a9",
X"26",
X"20",
X"24",
X"bc",
X"bd",
X"4c",
X"03",
X"bc",
X"4d",
X"03",
X"20",
X"33",
X"bd",
X"20",
X"af",
X"bc",
X"bd",
X"4e",
X"03",
X"4c",
X"31",
X"bd",
X"20",
X"a8",
X"bc",
X"20",
X"cd",
X"ab",
X"20",
X"af",
X"bc",
X"a5",
X"d4",
X"9d",
X"4c",
X"03",
X"a5",
X"d5",
X"9d",
X"4d",
X"03",
X"20",
X"cd",
X"ab",
X"20",
X"af",
X"bc",
X"a5",
X"d4",
X"9d",
X"4e",
X"03",
X"a9",
X"25",
X"85",
X"c0",
X"d0",
X"b1",
X"20",
X"a8",
X"bc",
X"20",
X"d7",
X"ab",
X"a5",
X"d4",
X"a6",
X"c1",
X"4c",
X"9b",
X"ba",
X"20",
X"51",
X"da",
X"20",
X"a8",
X"bc",
X"a9",
X"07",
X"85",
X"c0",
X"a0",
X"01",
X"20",
X"15",
X"bd",
X"20",
X"bb",
X"bc",
X"a0",
X"00",
X"b1",
X"f3",
X"4c",
X"31",
X"bd",
X"20",
X"0c",
X"ba",
X"a2",
X"06",
X"20",
X"c0",
X"ba",
X"d0",
X"e3",
X"20",
X"07",
X"bd",
X"85",
X"c1",
X"f0",
X"09",
X"a5",
X"c1",
X"0a",
X"0a",
X"0a",
X"0a",
X"aa",
X"10",
X"4e",
X"20",
X"0c",
X"b9",
X"20",
X"00",
X"bd",
X"10",
X"46",
X"a0",
X"00",
X"8c",
X"fe",
X"02",
X"c9",
X"80",
X"d0",
X"09",
X"84",
X"11",
X"a5",
X"ca",
X"f0",
X"37",
X"4c",
X"00",
X"a0",
X"a4",
X"c1",
X"c9",
X"88",
X"f0",
X"0f",
X"85",
X"b9",
X"c0",
X"07",
X"d0",
X"03",
X"20",
X"f7",
X"bc",
X"20",
X"5b",
X"bd",
X"4c",
X"34",
X"b9",
X"c0",
X"07",
X"d0",
X"ed",
X"a2",
X"5d",
X"e4",
X"c2",
X"d0",
X"e7",
X"20",
X"f7",
X"bc",
X"4c",
X"53",
X"a0",
X"20",
X"af",
X"bc",
X"f0",
X"0a",
X"a9",
X"0c",
X"d0",
X"2b",
X"20",
X"af",
X"bc",
X"bd",
X"43",
X"03",
X"60",
X"e6",
X"a8",
X"20",
X"cd",
X"ab",
X"a5",
X"d4",
X"60",
X"a0",
X"ff",
X"d0",
X"02",
X"a0",
X"00",
X"a9",
X"00",
X"9d",
X"49",
X"03",
X"98",
X"9d",
X"48",
X"03",
X"a5",
X"f4",
X"a4",
X"f3",
X"9d",
X"45",
X"03",
X"98",
X"9d",
X"44",
X"03",
X"a5",
X"c0",
X"9d",
X"42",
X"03",
X"4c",
X"56",
X"e4",
X"a0",
X"00",
X"48",
X"98",
X"48",
X"20",
X"06",
X"ac",
X"68",
X"85",
X"d5",
X"68",
X"85",
X"d4",
X"20",
X"aa",
X"d9",
X"4c",
X"0c",
X"ac",
X"a9",
X"00",
X"a2",
X"07",
X"9d",
X"00",
X"d2",
X"ca",
X"d0",
X"fa",
X"a0",
X"07",
X"84",
X"c1",
X"20",
X"f7",
X"bc",
X"c6",
X"c1",
X"d0",
X"f9",
X"60",
X"a9",
X"00",
X"85",
X"b4",
X"85",
X"b5",
X"60",
X"a2",
X"06",
X"86",
X"f2",
X"bd",
X"72",
X"bd",
X"20",
X"99",
X"ba",
X"a6",
X"f2",
X"ca",
X"10",
X"f3",
X"60",
X"9b",
X"59",
X"44",
X"41",
X"45",
X"52",
X"9b",
X"a2",
X"00",
X"f0",
X"e7",
X"20",
X"90",
X"ab",
X"a5",
X"d4",
X"85",
X"f3",
X"a5",
X"d5",
X"85",
X"f4",
X"a4",
X"d6",
X"a6",
X"d7",
X"f0",
X"02",
X"a0",
X"ff",
X"b1",
X"f3",
X"85",
X"97",
X"84",
X"98",
X"a9",
X"9b",
X"91",
X"f3",
X"85",
X"92",
X"60",
X"a4",
X"98",
X"a5",
X"97",
X"91",
X"f3",
X"a9",
X"00",
X"85",
X"92",
X"60",
X"20",
X"3e",
X"b8",
X"b0",
X"1b",
X"d0",
X"f9",
X"20",
X"cb",
X"bd",
X"c9",
X"0c",
X"f0",
X"24",
X"c9",
X"1e",
X"f0",
X"20",
X"c9",
X"04",
X"f0",
X"1c",
X"c9",
X"22",
X"f0",
X"18",
X"20",
X"f0",
X"b6",
X"20",
X"16",
X"b9",
X"20",
X"14",
X"b9",
X"20",
X"16",
X"b8",
X"b0",
X"f2",
X"a4",
X"b2",
X"88",
X"b1",
X"8a",
X"85",
X"a7",
X"c8",
X"b1",
X"8a",
X"60",
X"a6",
X"b4",
X"d0",
X"0e",
X"a9",
X"9b",
X"20",
X"99",
X"ba",
X"a6",
X"b4",
X"d0",
X"05",
X"a5",
X"c2",
X"20",
X"99",
X"ba",
X"a6",
X"b4",
X"a9",
X"05",
X"20",
X"be",
X"ba",
X"20",
X"0f",
X"bd",
X"4c",
X"bb",
X"bc",
X"20",
X"fd",
X"ab",
X"20",
X"26",
X"ad",
X"4c",
X"b2",
X"ab",
X"38",
X"60",
X"a9",
X"04",
X"24",
X"d4",
X"10",
X"06",
X"a9",
X"02",
X"d0",
X"02",
X"a9",
X"01",
X"85",
X"f0",
X"a5",
X"d4",
X"29",
X"7f",
X"85",
X"d4",
X"a9",
X"bd",
X"18",
X"65",
X"fb",
X"aa",
X"a0",
X"be",
X"20",
X"98",
X"dd",
X"20",
X"28",
X"db",
X"90",
X"01",
X"60",
X"a5",
X"d4",
X"29",
X"7f",
X"38",
X"e9",
X"40",
X"30",
X"2b",
X"c9",
X"04",
X"10",
X"cc",
X"aa",
X"b5",
X"d5",
X"85",
X"f1",
X"29",
X"10",
X"f0",
X"02",
X"a9",
X"02",
X"18",
X"65",
X"f1",
X"29",
X"03",
X"65",
X"f0",
X"85",
X"f0",
X"86",
X"f1",
X"20",
X"b6",
X"dd",
X"a6",
X"f1",
X"a9",
X"00",
X"95",
X"e2",
X"e8",
X"e0",
X"03",
X"90",
X"f9",
X"20",
X"60",
X"da",
X"46",
X"f0",
X"90",
X"0d",
X"20",
X"b6",
X"dd",
X"a2",
X"cf",
X"a0",
X"be",
X"20",
X"89",
X"dd",
X"20",
X"60",
X"da",
X"a2",
X"e6",
X"a0",
X"05",
X"20",
X"a7",
X"dd",
X"20",
X"b6",
X"dd",
X"20",
X"db",
X"da",
X"b0",
X"85",
X"a9",
X"06",
X"a2",
X"9f",
X"a0",
X"be",
X"20",
X"40",
X"dd",
X"a2",
X"e6",
X"a0",
X"05",
X"20",
X"98",
X"dd",
X"20",
X"db",
X"da",
X"46",
X"f0",
X"90",
X"09",
X"18",
X"a5",
X"d4",
X"f0",
X"04",
X"49",
X"80",
X"85",
X"d4",
X"60",
X"bd",
X"03",
X"55",
X"14",
X"99",
X"39",
X"3e",
X"01",
X"60",
X"44",
X"27",
X"52",
X"be",
X"46",
X"81",
X"75",
X"43",
X"55",
X"3f",
X"07",
X"96",
X"92",
X"62",
X"39",
X"bf",
X"64",
X"59",
X"64",
X"08",
X"67",
X"40",
X"01",
X"57",
X"07",
X"96",
X"32",
X"40",
X"90",
X"00",
X"00",
X"00",
X"00",
X"3f",
X"01",
X"74",
X"53",
X"29",
X"25",
X"40",
X"01",
X"00",
X"00",
X"00",
X"00",
X"a9",
X"00",
X"85",
X"f0",
X"85",
X"f1",
X"a5",
X"d4",
X"29",
X"7f",
X"c9",
X"40",
X"30",
X"15",
X"a5",
X"d4",
X"29",
X"80",
X"85",
X"f0",
X"e6",
X"f1",
X"a9",
X"7f",
X"25",
X"d4",
X"85",
X"d4",
X"a2",
X"ea",
X"a0",
X"df",
X"20",
X"95",
X"de",
X"a2",
X"e6",
X"a0",
X"05",
X"20",
X"a7",
X"dd",
X"20",
X"b6",
X"dd",
X"20",
X"db",
X"da",
X"b0",
X"39",
X"a9",
X"0b",
X"a2",
X"ae",
X"a0",
X"df",
X"20",
X"40",
X"dd",
X"b0",
X"2e",
X"a2",
X"e6",
X"a0",
X"05",
X"20",
X"98",
X"dd",
X"20",
X"db",
X"da",
X"b0",
X"22",
X"a5",
X"f1",
X"f0",
X"10",
X"a2",
X"f0",
X"a0",
X"df",
X"20",
X"98",
X"dd",
X"20",
X"66",
X"da",
X"a5",
X"f0",
X"05",
X"d4",
X"85",
X"d4",
X"a5",
X"fb",
X"f0",
X"0a",
X"a2",
X"c9",
X"a0",
X"be",
X"20",
X"98",
X"dd",
X"20",
X"28",
X"db",
X"60",
X"38",
X"60",
X"a9",
X"00",
X"85",
X"f1",
X"a5",
X"d4",
X"30",
X"f6",
X"c9",
X"3f",
X"f0",
X"17",
X"18",
X"69",
X"01",
X"85",
X"f1",
X"85",
X"e0",
X"a9",
X"01",
X"85",
X"e1",
X"a2",
X"04",
X"a9",
X"00",
X"95",
X"e2",
X"ca",
X"10",
X"fb",
X"20",
X"28",
X"db",
X"a9",
X"06",
X"85",
X"ef",
X"a2",
X"e6",
X"a0",
X"05",
X"20",
X"a7",
X"dd",
X"20",
X"b6",
X"dd",
X"a2",
X"f1",
X"a0",
X"ba",
X"20",
X"89",
X"dd",
X"20",
X"60",
X"da",
X"a2",
X"e6",
X"a0",
X"05",
X"20",
X"98",
X"dd",
X"20",
X"db",
X"da",
X"a2",
X"ec",
X"a0",
X"05",
X"20",
X"a7",
X"dd",
X"20",
X"b6",
X"dd",
X"a2",
X"e6",
X"a0",
X"05",
X"20",
X"89",
X"dd",
X"20",
X"28",
X"db",
X"a2",
X"ec",
X"a0",
X"05",
X"20",
X"98",
X"dd",
X"20",
X"60",
X"da",
X"a2",
X"6c",
X"a0",
X"df",
X"20",
X"98",
X"dd",
X"20",
X"db",
X"da",
X"a5",
X"d4",
X"f0",
X"0e",
X"a2",
X"ec",
X"a0",
X"05",
X"20",
X"98",
X"dd",
X"20",
X"66",
X"da",
X"c6",
X"ef",
X"10",
X"c6",
X"a2",
X"ec",
X"a0",
X"05",
X"20",
X"89",
X"dd",
X"a5",
X"f1",
X"f0",
X"23",
X"38",
X"e9",
X"40",
X"18",
X"6a",
X"18",
X"69",
X"40",
X"29",
X"7f",
X"85",
X"e0",
X"a5",
X"f1",
X"6a",
X"a9",
X"01",
X"90",
X"02",
X"a9",
X"10",
X"85",
X"e1",
X"a2",
X"04",
X"a9",
X"00",
X"95",
X"e2",
X"ca",
X"10",
X"fb",
X"20",
X"db",
X"da",
X"60",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"a0",
X"00",
X"05",
X"f0",
X"bf"

);
        signal rdata:std_logic_vector(7 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
			if we='1' then
				ROM(conv_integer(address)) <= data;
			end if;
                	q<=rdata;
                end if;
        end process;
end syn;
